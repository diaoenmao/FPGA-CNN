`define WIDTH 9
`define COUNTER_WIDTH 8
module sixteenbysixteen (
A1, A2, A3, A4, A5, A6, A7, A8, A9,
    
B1, B2, B3, B4, B5, B6, B7, B8, B9,
    
U1_in, U2_in, U3_in, U4_in, U5_in, U6_in, U7_in, U8_in, U9_in, U10_in, U11_in, U12_in, U13_in, U14_in, U15_in, U16_in,
U17_in, U18_in, U19_in, U20_in, U21_in, U22_in, U23_in, U24_in, U25_in, U26_in, U27_in, U28_in, U29_in, U30_in, U31_in, U32_in,
U33_in, U34_in, U35_in, U36_in, U37_in, U38_in, U39_in, U40_in, U41_in, U42_in, U43_in, U44_in, U45_in, U46_in, U47_in, U48_in,
U49_in, U50_in, U51_in, U52_in, U53_in, U54_in, U55_in, U56_in, U57_in, U58_in, U59_in, U60_in, U61_in, U62_in, U63_in, U64_in,
U65_in, U66_in, U67_in, U68_in, U69_in, U70_in, U71_in, U72_in, U73_in, U74_in, U75_in, U76_in, U77_in, U78_in, U79_in, U80_in,
U81_in, U82_in, U83_in, U84_in, U85_in, U86_in, U87_in, U88_in, U89_in, U90_in, U91_in, U92_in, U93_in, U94_in, U95_in, U96_in,
U97_in, U98_in, U99_in, U100_in, U101_in, U102_in, U103_in, U104_in, U105_in, U106_in, U107_in, U108_in, U109_in, U110_in, U111_in, U112_in,
U113_in, U114_in, U115_in, U116_in, U117_in, U118_in, U119_in, U120_in, U121_in, U122_in, U123_in, U124_in, U125_in, U126_in, U127_in, U128_in,

U129_in, U130_in, U131_in, U132_in, U133_in, U134_in, U135_in, U136_in, U137_in, U138_in, U139_in, U140_in, U141_in, U142_in, U143_in, U144_in,
U145_in, U146_in, U147_in, U148_in, U149_in, U150_in, U151_in, U152_in, U153_in, U154_in, U155_in, U156_in, U157_in, U158_in, U159_in, U160_in,
U161_in, U162_in, U163_in, U164_in, U165_in, U166_in, U167_in, U168_in, U169_in, U170_in, U171_in, U172_in, U173_in, U174_in, U175_in, U176_in,
U177_in, U178_in, U179_in, U180_in, U181_in, U182_in, U183_in, U184_in, U185_in, U186_in, U187_in, U188_in, U189_in, U190_in, U191_in, U192_in,
U193_in, U194_in, U195_in, U196_in, U197_in, U198_in, U199_in, U200_in, U201_in, U202_in, U203_in, U204_in, U205_in, U206_in, U207_in, U208_in,
U209_in, U210_in, U211_in, U212_in, U213_in, U214_in, U215_in, U216_in, U217_in, U218_in, U219_in, U220_in, U221_in, U222_in, U223_in, U224_in,
U225_in, U226_in, U227_in, U228_in, U229_in, U230_in, U231_in, U232_in, U233_in, U234_in, U235_in, U236_in, U237_in, U238_in, U239_in, U240_in,
U241_in, U242_in, U243_in, U244_in, U245_in, U246_in, U247_in, U248_in, U249_in, U250_in, U251_in, U252_in, U253_in, U254_in, U255_in, U256_in,
	
I,

Initial_X_in,

clk,

Y1_out, Y2_out, Y3_out, Y4_out, Y5_out, Y6_out, Y7_out, Y8_out, Y9_out, Y10_out, Y11_out, Y12_out, Y13_out, Y14_out, Y15_out, Y16_out,
Y17_out, Y18_out, Y19_out, Y20_out, Y21_out, Y22_out, Y23_out, Y24_out, Y25_out, Y26_out, Y27_out, Y28_out, Y29_out, Y30_out, Y31_out, Y32_out,
Y33_out, Y34_out, Y35_out, Y36_out, Y37_out, Y38_out, Y39_out, Y40_out, Y41_out, Y42_out, Y43_out, Y44_out, Y45_out, Y46_out, Y47_out, Y48_out,
Y49_out, Y50_out, Y51_out, Y52_out, Y53_out, Y54_out, Y55_out, Y56_out, Y57_out, Y58_out, Y59_out, Y60_out, Y61_out, Y62_out, Y63_out, Y64_out,
Y65_out, Y66_out, Y67_out, Y68_out, Y69_out, Y70_out, Y71_out, Y72_out, Y73_out, Y74_out, Y75_out, Y76_out, Y77_out, Y78_out, Y79_out, Y80_out,
Y81_out, Y82_out, Y83_out, Y84_out, Y85_out, Y86_out, Y87_out, Y88_out, Y89_out, Y90_out, Y91_out, Y92_out, Y93_out, Y94_out, Y95_out, Y96_out,
Y97_out, Y98_out, Y99_out, Y100_out, Y101_out, Y102_out, Y103_out, Y104_out, Y105_out, Y106_out, Y107_out, Y108_out, Y109_out, Y110_out, Y111_out, Y112_out,
Y113_out, Y114_out, Y115_out, Y116_out, Y117_out, Y118_out, Y119_out, Y120_out, Y121_out, Y122_out, Y123_out, Y124_out, Y125_out, Y126_out, Y127_out, Y128_out,

Y129_out, Y130_out, Y131_out, Y132_out, Y133_out, Y134_out, Y135_out, Y136_out, Y137_out, Y138_out, Y139_out, Y140_out, Y141_out, Y142_out, Y143_out, Y144_out,
Y145_out, Y146_out, Y147_out, Y148_out, Y149_out, Y150_out, Y151_out, Y152_out, Y153_out, Y154_out, Y155_out, Y156_out, Y157_out, Y158_out, Y159_out, Y160_out,
Y161_out, Y162_out, Y163_out, Y164_out, Y165_out, Y166_out, Y167_out, Y168_out, Y169_out, Y170_out, Y171_out, Y172_out, Y173_out, Y174_out, Y175_out, Y176_out,
Y177_out, Y178_out, Y179_out, Y180_out, Y181_out, Y182_out, Y183_out, Y184_out, Y185_out, Y186_out, Y187_out, Y188_out, Y189_out, Y190_out, Y191_out, Y192_out,
Y193_out, Y194_out, Y195_out, Y196_out, Y197_out, Y198_out, Y199_out, Y200_out, Y201_out, Y202_out, Y203_out, Y204_out, Y205_out, Y206_out, Y207_out, Y208_out,
Y209_out, Y210_out, Y211_out, Y212_out, Y213_out, Y214_out, Y215_out, Y216_out, Y217_out, Y218_out, Y219_out, Y220_out, Y221_out, Y222_out, Y223_out, Y224_out,
Y225_out, Y226_out, Y227_out, Y228_out, Y229_out, Y230_out, Y231_out, Y232_out, Y233_out, Y234_out, Y235_out, Y236_out, Y237_out, Y238_out, Y239_out, Y240_out,
Y241_out, Y242_out, Y243_out, Y244_out, Y245_out, Y246_out, Y247_out, Y248_out, Y249_out, Y250_out, Y251_out, Y252_out, Y253_out, Y254_out, Y255_out, Y256_out

  );
	input wire clk;
	input wire signed [`WIDTH - 1:0] A1, A2, A3, A4, A5, A6, A7, A8, A9;
	input wire signed [`WIDTH - 1:0] B1, B2, B3, B4, B5, B6, B7, B8, B9;
	input wire signed [`WIDTH - 1:0] U1_in, U2_in, U3_in, U4_in, U5_in, U6_in, U7_in, U8_in, U9_in, U10_in, U11_in, U12_in, U13_in, U14_in, U15_in, U16_in;
	input wire signed [`WIDTH - 1:0] U17_in, U18_in, U19_in, U20_in, U21_in, U22_in, U23_in, U24_in, U25_in, U26_in, U27_in, U28_in, U29_in, U30_in, U31_in, U32_in;
	input wire signed [`WIDTH - 1:0] U33_in, U34_in, U35_in, U36_in, U37_in, U38_in, U39_in, U40_in, U41_in, U42_in, U43_in, U44_in, U45_in, U46_in, U47_in, U48_in;
	input wire signed [`WIDTH - 1:0] U49_in, U50_in, U51_in, U52_in, U53_in, U54_in, U55_in, U56_in, U57_in, U58_in, U59_in, U60_in, U61_in, U62_in, U63_in, U64_in;
	input wire signed [`WIDTH - 1:0] U65_in, U66_in, U67_in, U68_in, U69_in, U70_in, U71_in, U72_in, U73_in, U74_in, U75_in, U76_in, U77_in, U78_in, U79_in, U80_in;
	input wire signed [`WIDTH - 1:0] U81_in, U82_in, U83_in, U84_in, U85_in, U86_in, U87_in, U88_in, U89_in, U90_in, U91_in, U92_in, U93_in, U94_in, U95_in, U96_in;
	input wire signed [`WIDTH - 1:0] U97_in, U98_in, U99_in, U100_in, U101_in, U102_in, U103_in, U104_in, U105_in, U106_in, U107_in, U108_in, U109_in, U110_in, U111_in, U112_in;
	input wire signed [`WIDTH - 1:0] U113_in, U114_in, U115_in, U116_in, U117_in, U118_in, U119_in, U120_in, U121_in, U122_in, U123_in, U124_in, U125_in, U126_in, U127_in, U128_in;

	input wire signed [`WIDTH - 1:0] U129_in, U130_in, U131_in, U132_in, U133_in, U134_in, U135_in, U136_in, U137_in, U138_in, U139_in, U140_in, U141_in, U142_in, U143_in, U144_in;
	input wire signed [`WIDTH - 1:0] U145_in, U146_in, U147_in, U148_in, U149_in, U150_in, U151_in, U152_in, U153_in, U154_in, U155_in, U156_in, U157_in, U158_in, U159_in, U160_in;
	input wire signed [`WIDTH - 1:0] U161_in, U162_in, U163_in, U164_in, U165_in, U166_in, U167_in, U168_in, U169_in, U170_in, U171_in, U172_in, U173_in, U174_in, U175_in, U176_in;
	input wire signed [`WIDTH - 1:0] U177_in, U178_in, U179_in, U180_in, U181_in, U182_in, U183_in, U184_in, U185_in, U186_in, U187_in, U188_in, U189_in, U190_in, U191_in, U192_in;
	input wire signed [`WIDTH - 1:0] U193_in, U194_in, U195_in, U196_in, U197_in, U198_in, U199_in, U200_in, U201_in, U202_in, U203_in, U204_in, U205_in, U206_in, U207_in, U208_in;
	input wire signed [`WIDTH - 1:0] U209_in, U210_in, U211_in, U212_in, U213_in, U214_in, U215_in, U216_in, U217_in, U218_in, U219_in, U220_in, U221_in, U222_in, U223_in, U224_in;
	input wire signed [`WIDTH - 1:0] U225_in, U226_in, U227_in, U228_in, U229_in, U230_in, U231_in, U232_in, U233_in, U234_in, U235_in, U236_in, U237_in, U238_in, U239_in, U240_in;
	input wire signed [`WIDTH - 1:0] U241_in, U242_in, U243_in, U244_in, U245_in, U246_in, U247_in, U248_in, U249_in, U250_in, U251_in, U252_in, U253_in, U254_in, U255_in, U256_in;
	
	input wire signed [`WIDTH - 1:0] I;
	input wire signed [2 * `WIDTH - 1:0] Initial_X_in;
	reg signed [2 * `WIDTH - 1:0] Initial_X;
	reg signed [`WIDTH - 1:0] U1, U2, U3, U4, U5, U6, U7, U8, U9;
	reg signed [2 * `WIDTH - 1:0] Y1_in = `WIDTH'b0, Y2_in = `WIDTH'b0, Y3_in = `WIDTH'b0, Y4_in = `WIDTH'b0, Y5_in = `WIDTH'b0, Y6_in = `WIDTH'b0, Y7_in = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y8_in = `WIDTH'b0, Y9_in = `WIDTH'b0, Y10_in = `WIDTH'b0, Y11_in = `WIDTH'b0, Y12_in = `WIDTH'b0, Y13_in = `WIDTH'b0, Y14_in = `WIDTH'b0, Y15_in = `WIDTH'b0, Y16_in = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y1, Y2 , Y3, Y4, Y5, Y6, Y7, Y8, Y9;
	reg [`COUNTER_WIDTH - 1:0] counter = `COUNTER_WIDTH'b0;
	wire signed [2 * `WIDTH - 1:0] onebyoneout;
	
	reg signed [2 * `WIDTH - 1:0] Y1_next = `WIDTH'b0, Y2_next = `WIDTH'b0, Y3_next = `WIDTH'b0, Y4_next = `WIDTH'b0, Y5_next = `WIDTH'b0, Y6_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y7_next = `WIDTH'b0, Y8_next = `WIDTH'b0, Y9_next = `WIDTH'b0, Y10_next = `WIDTH'b0, Y11_next = `WIDTH'b0, Y12_next = `WIDTH'b0, Y13_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y14_next = `WIDTH'b0, Y15_next = `WIDTH'b0, Y16_next = `WIDTH'b0, Y17_next = `WIDTH'b0, Y18_next = `WIDTH'b0, Y19_next = `WIDTH'b0, Y20_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y21_next = `WIDTH'b0, Y22_next = `WIDTH'b0, Y23_next = `WIDTH'b0, Y24_next = `WIDTH'b0, Y25_next = `WIDTH'b0, Y26_next = `WIDTH'b0, Y27_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y28_next = `WIDTH'b0, Y29_next = `WIDTH'b0, Y30_next = `WIDTH'b0, Y31_next = `WIDTH'b0, Y32_next = `WIDTH'b0, Y33_next = `WIDTH'b0, Y34_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y35_next = `WIDTH'b0, Y36_next = `WIDTH'b0, Y37_next = `WIDTH'b0, Y38_next = `WIDTH'b0, Y39_next = `WIDTH'b0, Y40_next = `WIDTH'b0, Y41_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y42_next = `WIDTH'b0, Y43_next = `WIDTH'b0, Y44_next = `WIDTH'b0, Y45_next = `WIDTH'b0, Y46_next = `WIDTH'b0, Y47_next = `WIDTH'b0, Y48_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y49_next = `WIDTH'b0, Y50_next = `WIDTH'b0, Y51_next = `WIDTH'b0, Y52_next = `WIDTH'b0, Y53_next = `WIDTH'b0, Y54_next = `WIDTH'b0, Y55_next = `WIDTH'b0; 
	reg signed [2 * `WIDTH - 1:0] Y56_next = `WIDTH'b0, Y57_next = `WIDTH'b0, Y58_next = `WIDTH'b0, Y59_next = `WIDTH'b0, Y60_next = `WIDTH'b0, Y61_next = `WIDTH'b0, Y62_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y63_next = `WIDTH'b0, Y64_next = `WIDTH'b0, Y65_next = `WIDTH'b0, Y66_next = `WIDTH'b0, Y67_next = `WIDTH'b0, Y68_next = `WIDTH'b0, Y69_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y70_next = `WIDTH'b0, Y71_next = `WIDTH'b0, Y72_next = `WIDTH'b0, Y73_next = `WIDTH'b0, Y74_next = `WIDTH'b0, Y75_next = `WIDTH'b0, Y76_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y77_next = `WIDTH'b0, Y78_next = `WIDTH'b0, Y79_next = `WIDTH'b0, Y80_next = `WIDTH'b0, Y81_next = `WIDTH'b0, Y82_next = `WIDTH'b0, Y83_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y84_next = `WIDTH'b0, Y85_next = `WIDTH'b0, Y86_next = `WIDTH'b0, Y87_next = `WIDTH'b0, Y88_next = `WIDTH'b0, Y89_next = `WIDTH'b0, Y90_next = `WIDTH'b0; 
	reg signed [2 * `WIDTH - 1:0] Y91_next = `WIDTH'b0, Y92_next = `WIDTH'b0, Y93_next = `WIDTH'b0, Y94_next = `WIDTH'b0, Y95_next = `WIDTH'b0, Y96_next = `WIDTH'b0, Y97_next = `WIDTH'b0; 
	reg signed [2 * `WIDTH - 1:0] Y98_next = `WIDTH'b0, Y99_next = `WIDTH'b0, Y100_next = `WIDTH'b0, Y101_next = `WIDTH'b0, Y102_next = `WIDTH'b0, Y103_next = `WIDTH'b0, Y104_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y105_next = `WIDTH'b0, Y106_next = `WIDTH'b0, Y107_next = `WIDTH'b0, Y108_next = `WIDTH'b0, Y109_next = `WIDTH'b0, Y110_next = `WIDTH'b0, Y111_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y112_next = `WIDTH'b0, Y113_next = `WIDTH'b0, Y114_next = `WIDTH'b0, Y115_next = `WIDTH'b0, Y116_next = `WIDTH'b0, Y117_next = `WIDTH'b0, Y118_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y119_next = `WIDTH'b0, Y120_next = `WIDTH'b0, Y121_next = `WIDTH'b0, Y122_next = `WIDTH'b0, Y123_next = `WIDTH'b0, Y124_next = `WIDTH'b0, Y125_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y126_next = `WIDTH'b0, Y127_next = `WIDTH'b0, Y128_next = `WIDTH'b0, Y129_next = `WIDTH'b0, Y130_next = `WIDTH'b0, Y131_next = `WIDTH'b0, Y132_next = `WIDTH'b0;	
	reg signed [2 * `WIDTH - 1:0] Y133_next = `WIDTH'b0, Y134_next = `WIDTH'b0, Y135_next = `WIDTH'b0, Y136_next = `WIDTH'b0, Y137_next = `WIDTH'b0, Y138_next = `WIDTH'b0, Y139_next = `WIDTH'b0;	
	reg signed [2 * `WIDTH - 1:0] Y140_next = `WIDTH'b0, Y141_next = `WIDTH'b0, Y142_next = `WIDTH'b0, Y143_next = `WIDTH'b0, Y144_next = `WIDTH'b0, Y145_next = `WIDTH'b0, Y146_next = `WIDTH'b0;	
	reg signed [2 * `WIDTH - 1:0] Y147_next = `WIDTH'b0, Y148_next = `WIDTH'b0, Y149_next = `WIDTH'b0, Y150_next = `WIDTH'b0, Y151_next = `WIDTH'b0, Y152_next = `WIDTH'b0, Y153_next = `WIDTH'b0;	
	reg signed [2 * `WIDTH - 1:0] Y154_next = `WIDTH'b0, Y155_next = `WIDTH'b0, Y156_next = `WIDTH'b0, Y157_next = `WIDTH'b0, Y158_next = `WIDTH'b0, Y159_next = `WIDTH'b0, Y160_next = `WIDTH'b0; 	
	reg signed [2 * `WIDTH - 1:0] Y161_next = `WIDTH'b0, Y162_next = `WIDTH'b0, Y163_next = `WIDTH'b0, Y164_next = `WIDTH'b0, Y165_next = `WIDTH'b0, Y166_next = `WIDTH'b0, Y167_next = `WIDTH'b0; 
	reg signed [2 * `WIDTH - 1:0] Y168_next = `WIDTH'b0, Y169_next = `WIDTH'b0, Y170_next = `WIDTH'b0, Y171_next = `WIDTH'b0, Y172_next = `WIDTH'b0, Y173_next = `WIDTH'b0, Y174_next = `WIDTH'b0;	
	reg signed [2 * `WIDTH - 1:0] Y175_next = `WIDTH'b0, Y176_next = `WIDTH'b0, Y177_next = `WIDTH'b0, Y178_next = `WIDTH'b0, Y179_next = `WIDTH'b0, Y180_next = `WIDTH'b0, Y181_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y182_next = `WIDTH'b0, Y183_next = `WIDTH'b0, Y184_next = `WIDTH'b0, Y185_next = `WIDTH'b0, Y186_next = `WIDTH'b0, Y187_next = `WIDTH'b0, Y188_next = `WIDTH'b0; 	
	reg signed [2 * `WIDTH - 1:0] Y189_next = `WIDTH'b0, Y190_next = `WIDTH'b0, Y191_next = `WIDTH'b0, Y192_next = `WIDTH'b0, Y193_next = `WIDTH'b0, Y194_next = `WIDTH'b0, Y195_next = `WIDTH'b0;	
	reg signed [2 * `WIDTH - 1:0] Y196_next = `WIDTH'b0, Y197_next = `WIDTH'b0, Y198_next = `WIDTH'b0, Y199_next = `WIDTH'b0, Y200_next = `WIDTH'b0, Y201_next = `WIDTH'b0, Y202_next = `WIDTH'b0;	
	reg signed [2 * `WIDTH - 1:0] Y203_next = `WIDTH'b0, Y204_next = `WIDTH'b0, Y205_next = `WIDTH'b0, Y206_next = `WIDTH'b0, Y207_next = `WIDTH'b0, Y208_next = `WIDTH'b0, Y209_next = `WIDTH'b0;	
	reg signed [2 * `WIDTH - 1:0] Y210_next = `WIDTH'b0, Y211_next = `WIDTH'b0, Y212_next = `WIDTH'b0, Y213_next = `WIDTH'b0, Y214_next = `WIDTH'b0, Y215_next = `WIDTH'b0, Y216_next = `WIDTH'b0;	
	reg signed [2 * `WIDTH - 1:0] Y217_next = `WIDTH'b0, Y218_next = `WIDTH'b0, Y219_next = `WIDTH'b0, Y220_next = `WIDTH'b0, Y221_next = `WIDTH'b0, Y222_next = `WIDTH'b0, Y223_next = `WIDTH'b0;	
	reg signed [2 * `WIDTH - 1:0] Y224_next = `WIDTH'b0, Y225_next = `WIDTH'b0, Y226_next = `WIDTH'b0, Y227_next = `WIDTH'b0, Y228_next = `WIDTH'b0, Y229_next = `WIDTH'b0, Y230_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y231_next = `WIDTH'b0, Y232_next = `WIDTH'b0, Y233_next = `WIDTH'b0, Y234_next = `WIDTH'b0, Y235_next = `WIDTH'b0, Y236_next = `WIDTH'b0, Y237_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y238_next = `WIDTH'b0, Y239_next = `WIDTH'b0, Y240_next = `WIDTH'b0, Y241_next = `WIDTH'b0, Y242_next = `WIDTH'b0, Y243_next = `WIDTH'b0, Y244_next = `WIDTH'b0; 
	reg signed [2 * `WIDTH - 1:0] Y245_next = `WIDTH'b0, Y246_next = `WIDTH'b0, Y247_next = `WIDTH'b0, Y248_next = `WIDTH'b0, Y249_next = `WIDTH'b0, Y250_next = `WIDTH'b0, Y251_next = `WIDTH'b0;
	reg signed [2 * `WIDTH - 1:0] Y252_next = `WIDTH'b0, Y253_next = `WIDTH'b0, Y254_next = `WIDTH'b0, Y255_next = `WIDTH'b0, Y256_next = `WIDTH'b0;
	
						
	output wire signed [2 * `WIDTH - 1:0] Y1_out, Y2_out, Y3_out, Y4_out, Y5_out, Y6_out, Y7_out, Y8_out, Y9_out, Y10_out, Y11_out, Y12_out, Y13_out, Y14_out, Y15_out, Y16_out;
	output wire signed [2 * `WIDTH - 1:0] Y17_out, Y18_out, Y19_out, Y20_out, Y21_out, Y22_out, Y23_out, Y24_out, Y25_out, Y26_out, Y27_out, Y28_out, Y29_out, Y30_out, Y31_out, Y32_out,
	output wire signed [2 * `WIDTH - 1:0] Y33_out, Y34_out, Y35_out, Y36_out, Y37_out, Y38_out, Y39_out, Y40_out, Y41_out, Y42_out, Y43_out, Y44_out, Y45_out, Y46_out, Y47_out, Y48_out,
	output wire signed [2 * `WIDTH - 1:0] Y49_out, Y50_out, Y51_out, Y52_out, Y53_out, Y54_out, Y55_out, Y56_out, Y57_out, Y58_out, Y59_out, Y60_out, Y61_out, Y62_out, Y63_out, Y64_out,
	output wire signed [2 * `WIDTH - 1:0] Y65_out, Y66_out, Y67_out, Y68_out, Y69_out, Y70_out, Y71_out, Y72_out, Y73_out, Y74_out, Y75_out, Y76_out, Y77_out, Y78_out, Y79_out, Y80_out,
	output wire signed [2 * `WIDTH - 1:0] Y81_out, Y82_out, Y83_out, Y84_out, Y85_out, Y86_out, Y87_out, Y88_out, Y89_out, Y90_out, Y91_out, Y92_out, Y93_out, Y94_out, Y95_out, Y96_out,
	output wire signed [2 * `WIDTH - 1:0] Y97_out, Y98_out, Y99_out, Y100_out, Y101_out, Y102_out, Y103_out, Y104_out, Y105_out, Y106_out, Y107_out, Y108_out, Y109_out, Y110_out, Y111_out, Y112_out,
	output wire signed [2 * `WIDTH - 1:0] Y113_out, Y114_out, Y115_out, Y116_out, Y117_out, Y118_out, Y119_out, Y120_out, Y121_out, Y122_out, Y123_out, Y124_out, Y125_out, Y126_out, Y127_out, Y128_out,

	output wire signed [2 * `WIDTH - 1:0] Y129_out, Y130_out, Y131_out, Y132_out, Y133_out, Y134_out, Y135_out, Y136_out, Y137_out, Y138_out, Y139_out, Y140_out, Y141_out, Y142_out, Y143_out, Y144_out,
	output wire signed [2 * `WIDTH - 1:0] Y145_out, Y146_out, Y147_out, Y148_out, Y149_out, Y150_out, Y151_out, Y152_out, Y153_out, Y154_out, Y155_out, Y156_out, Y157_out, Y158_out, Y159_out, Y160_out,
	output wire signed [2 * `WIDTH - 1:0] Y161_out, Y162_out, Y163_out, Y164_out, Y165_out, Y166_out, Y167_out, Y168_out, Y169_out, Y170_out, Y171_out, Y172_out, Y173_out, Y174_out, Y175_out, Y176_out,
	output wire signed [2 * `WIDTH - 1:0] Y177_out, Y178_out, Y179_out, Y180_out, Y181_out, Y182_out, Y183_out, Y184_out, Y185_out, Y186_out, Y187_out, Y188_out, Y189_out, Y190_out, Y191_out, Y192_out,
	output wire signed [2 * `WIDTH - 1:0] Y193_out, Y194_out, Y195_out, Y196_out, Y197_out, Y198_out, Y199_out, Y200_out, Y201_out, Y202_out, Y203_out, Y204_out, Y205_out, Y206_out, Y207_out, Y208_out,
	output wire signed [2 * `WIDTH - 1:0] Y209_out, Y210_out, Y211_out, Y212_out, Y213_out, Y214_out, Y215_out, Y216_out, Y217_out, Y218_out, Y219_out, Y220_out, Y221_out, Y222_out, Y223_out, Y224_out,
	output wire signed [2 * `WIDTH - 1:0] Y225_out, Y226_out, Y227_out, Y228_out, Y229_out, Y230_out, Y231_out, Y232_out, Y233_out, Y234_out, Y235_out, Y236_out, Y237_out, Y238_out, Y239_out, Y240_out,
	output wire signed [2 * `WIDTH - 1:0] Y241_out, Y242_out, Y243_out, Y244_out, Y245_out, Y246_out, Y247_out, Y248_out, Y249_out, Y250_out, Y251_out, Y252_out, Y253_out, Y254_out, Y255_out, Y256_out
	
    reg initial_flag = 1'b1;
    
    
assign Y1_out = Y1_next;
assign Y2_out = Y2_next;
assign Y3_out = Y3_next;
assign Y4_out = Y4_next;
assign Y5_out = Y5_next;
assign Y6_out = Y6_next;
assign Y7_out = Y7_next;
assign Y8_out = Y8_next;
assign Y9_out = Y9_next;
assign Y10_out = Y10_next;
assign Y11_out = Y11_next;
assign Y12_out = Y12_next;
assign Y13_out = Y13_next;
assign Y14_out = Y14_next;
assign Y15_out = Y15_next;
assign Y16_out = Y16_next;
assign Y17_out = Y17_next;
assign Y18_out = Y18_next;
assign Y19_out = Y19_next;
assign Y20_out = Y20_next;
assign Y21_out = Y21_next;
assign Y22_out = Y22_next;
assign Y23_out = Y23_next;
assign Y24_out = Y24_next;
assign Y25_out = Y25_next;
assign Y26_out = Y26_next;
assign Y27_out = Y27_next;
assign Y28_out = Y28_next;
assign Y29_out = Y29_next;
assign Y30_out = Y30_next;
assign Y31_out = Y31_next;
assign Y32_out = Y32_next;
assign Y33_out = Y33_next;
assign Y34_out = Y34_next;
assign Y35_out = Y35_next;
assign Y36_out = Y36_next;
assign Y37_out = Y37_next;
assign Y38_out = Y38_next;
assign Y39_out = Y39_next;
assign Y40_out = Y40_next;
assign Y41_out = Y41_next;
assign Y42_out = Y42_next;
assign Y43_out = Y43_next;
assign Y44_out = Y44_next;
assign Y45_out = Y45_next;
assign Y46_out = Y46_next;
assign Y47_out = Y47_next;
assign Y48_out = Y48_next;
assign Y49_out = Y49_next;
assign Y50_out = Y50_next;
assign Y51_out = Y51_next;
assign Y52_out = Y52_next;
assign Y53_out = Y53_next;
assign Y54_out = Y54_next;
assign Y55_out = Y55_next;
assign Y56_out = Y56_next;
assign Y57_out = Y57_next;
assign Y58_out = Y58_next;
assign Y59_out = Y59_next;
assign Y60_out = Y60_next;
assign Y61_out = Y61_next;
assign Y62_out = Y62_next;
assign Y63_out = Y63_next;
assign Y64_out = Y64_next;
assign Y65_out = Y65_next;
assign Y66_out = Y66_next;
assign Y67_out = Y67_next;
assign Y68_out = Y68_next;
assign Y69_out = Y69_next;
assign Y70_out = Y70_next;
assign Y71_out = Y71_next;
assign Y72_out = Y72_next;
assign Y73_out = Y73_next;
assign Y74_out = Y74_next;
assign Y75_out = Y75_next;
assign Y76_out = Y76_next;
assign Y77_out = Y77_next;
assign Y78_out = Y78_next;
assign Y79_out = Y79_next;
assign Y80_out = Y80_next;
assign Y81_out = Y81_next;
assign Y82_out = Y82_next;
assign Y83_out = Y83_next;
assign Y84_out = Y84_next;
assign Y85_out = Y85_next;
assign Y86_out = Y86_next;
assign Y87_out = Y87_next;
assign Y88_out = Y88_next;
assign Y89_out = Y89_next;
assign Y90_out = Y90_next;
assign Y91_out = Y91_next;
assign Y92_out = Y92_next;
assign Y93_out = Y93_next;
assign Y94_out = Y94_next;
assign Y95_out = Y95_next;
assign Y96_out = Y96_next;
assign Y97_out = Y97_next;
assign Y98_out = Y98_next;
assign Y99_out = Y99_next;
assign Y100_out = Y100_next;
assign Y101_out = Y101_next;
assign Y102_out = Y102_next;
assign Y103_out = Y103_next;
assign Y104_out = Y104_next;
assign Y105_out = Y105_next;
assign Y106_out = Y106_next;
assign Y107_out = Y107_next;
assign Y108_out = Y108_next;
assign Y109_out = Y109_next;
assign Y110_out = Y110_next;
assign Y111_out = Y111_next;
assign Y112_out = Y112_next;
assign Y113_out = Y113_next;
assign Y114_out = Y114_next;
assign Y115_out = Y115_next;
assign Y116_out = Y116_next;
assign Y117_out = Y117_next;
assign Y118_out = Y118_next;
assign Y119_out = Y119_next;
assign Y120_out = Y120_next;
assign Y121_out = Y121_next;
assign Y122_out = Y122_next;
assign Y123_out = Y123_next;
assign Y124_out = Y124_next;
assign Y125_out = Y125_next;
assign Y126_out = Y126_next;
assign Y127_out = Y127_next;
assign Y128_out = Y128_next;
assign Y129_out = Y129_next;
assign Y130_out = Y130_next;
assign Y131_out = Y131_next;
assign Y132_out = Y132_next;
assign Y133_out = Y133_next;
assign Y134_out = Y134_next;
assign Y135_out = Y135_next;
assign Y136_out = Y136_next;
assign Y137_out = Y137_next;
assign Y138_out = Y138_next;
assign Y139_out = Y139_next;
assign Y140_out = Y140_next;
assign Y141_out = Y141_next;
assign Y142_out = Y142_next;
assign Y143_out = Y143_next;
assign Y144_out = Y144_next;
assign Y145_out = Y145_next;
assign Y146_out = Y146_next;
assign Y147_out = Y147_next;
assign Y148_out = Y148_next;
assign Y149_out = Y149_next;
assign Y150_out = Y150_next;
assign Y151_out = Y151_next;
assign Y152_out = Y152_next;
assign Y153_out = Y153_next;
assign Y154_out = Y154_next;
assign Y155_out = Y155_next;
assign Y156_out = Y156_next;
assign Y157_out = Y157_next;
assign Y158_out = Y158_next;
assign Y159_out = Y159_next;
assign Y160_out = Y160_next;
assign Y161_out = Y161_next;
assign Y162_out = Y162_next;
assign Y163_out = Y163_next;
assign Y164_out = Y164_next;
assign Y165_out = Y165_next;
assign Y166_out = Y166_next;
assign Y167_out = Y167_next;
assign Y168_out = Y168_next;
assign Y169_out = Y169_next;
assign Y170_out = Y170_next;
assign Y171_out = Y171_next;
assign Y172_out = Y172_next;
assign Y173_out = Y173_next;
assign Y174_out = Y174_next;
assign Y175_out = Y175_next;
assign Y176_out = Y176_next;
assign Y177_out = Y177_next;
assign Y178_out = Y178_next;
assign Y179_out = Y179_next;
assign Y180_out = Y180_next;
assign Y181_out = Y181_next;
assign Y182_out = Y182_next;
assign Y183_out = Y183_next;
assign Y184_out = Y184_next;
assign Y185_out = Y185_next;
assign Y186_out = Y186_next;
assign Y187_out = Y187_next;
assign Y188_out = Y188_next;
assign Y189_out = Y189_next;
assign Y190_out = Y190_next;
assign Y191_out = Y191_next;
assign Y192_out = Y192_next;
assign Y193_out = Y193_next;
assign Y194_out = Y194_next;
assign Y195_out = Y195_next;
assign Y196_out = Y196_next;
assign Y197_out = Y197_next;
assign Y198_out = Y198_next;
assign Y199_out = Y199_next;
assign Y200_out = Y200_next;
assign Y201_out = Y201_next;
assign Y202_out = Y202_next;
assign Y203_out = Y203_next;
assign Y204_out = Y204_next;
assign Y205_out = Y205_next;
assign Y206_out = Y206_next;
assign Y207_out = Y207_next;
assign Y208_out = Y208_next;
assign Y209_out = Y209_next;
assign Y210_out = Y210_next;
assign Y211_out = Y211_next;
assign Y212_out = Y212_next;
assign Y213_out = Y213_next;
assign Y214_out = Y214_next;
assign Y215_out = Y215_next;
assign Y216_out = Y216_next;
assign Y217_out = Y217_next;
assign Y218_out = Y218_next;
assign Y219_out = Y219_next;
assign Y220_out = Y220_next;
assign Y221_out = Y221_next;
assign Y222_out = Y222_next;
assign Y223_out = Y223_next;
assign Y224_out = Y224_next;
assign Y225_out = Y225_next;
assign Y226_out = Y226_next;
assign Y227_out = Y227_next;
assign Y228_out = Y228_next;
assign Y229_out = Y229_next;
assign Y230_out = Y230_next;
assign Y231_out = Y231_next;
assign Y232_out = Y232_next;
assign Y233_out = Y233_next;
assign Y234_out = Y234_next;
assign Y235_out = Y235_next;
assign Y236_out = Y236_next;
assign Y237_out = Y237_next;
assign Y238_out = Y238_next;
assign Y239_out = Y239_next;
assign Y240_out = Y240_next;
assign Y241_out = Y241_next;
assign Y242_out = Y242_next;
assign Y243_out = Y243_next;
assign Y244_out = Y244_next;
assign Y245_out = Y245_next;
assign Y246_out = Y246_next;
assign Y247_out = Y247_next;
assign Y248_out = Y248_next;
assign Y249_out = Y249_next;
assign Y250_out = Y250_next;
assign Y251_out = Y251_next;
assign Y252_out = Y252_next;
assign Y253_out = Y253_next;
assign Y254_out = Y254_next;
assign Y255_out = Y255_next;
assign Y256_out = Y256_next;






always  @ (posedge clk)
begin
  
  if (counter == `COUNTER_WIDTH'b0) begin // 1    
	
	if (initial_flag == 1'b0) begin
	    Initial_X = {(2 * `WIDTH){1'b0}};
	    
		Y256_next = onebyoneout;

		Y1_in = Y1_next;
		Y2_in = Y2_next;
		Y3_in = Y3_next;
		Y4_in = Y4_next;
		Y5_in = Y5_next;
		Y6_in = Y6_next;
		Y7_in = Y7_next;
		Y8_in = Y8_next;
		Y9_in = Y9_next;
		Y10_in = Y10_next;
		Y11_in = Y11_next;
		Y12_in = Y12_next;
		Y13_in = Y13_next;
		Y14_in = Y14_next;
		Y15_in = Y15_next;
		Y16_in = Y16_next;
		Y17_in = Y17_next;
		Y18_in = Y18_next;
		Y19_in = Y19_next;
		Y20_in = Y20_next;
		Y21_in = Y21_next;
		Y22_in = Y22_next;
		Y23_in = Y23_next;
		Y24_in = Y24_next;
		Y25_in = Y25_next;
		Y26_in = Y26_next;
		Y27_in = Y27_next;
		Y28_in = Y28_next;
		Y29_in = Y29_next;
		Y30_in = Y30_next;
		Y31_in = Y31_next;
		Y32_in = Y32_next;
		Y33_in = Y33_next;
		Y34_in = Y34_next;
		Y35_in = Y35_next;
		Y36_in = Y36_next;
		Y37_in = Y37_next;
		Y38_in = Y38_next;
		Y39_in = Y39_next;
		Y40_in = Y40_next;
		Y41_in = Y41_next;
		Y42_in = Y42_next;
		Y43_in = Y43_next;
		Y44_in = Y44_next;
		Y45_in = Y45_next;
		Y46_in = Y46_next;
		Y47_in = Y47_next;
		Y48_in = Y48_next;
		Y49_in = Y49_next;
		Y50_in = Y50_next;
		Y51_in = Y51_next;
		Y52_in = Y52_next;
		Y53_in = Y53_next;
		Y54_in = Y54_next;
		Y55_in = Y55_next;
		Y56_in = Y56_next;
		Y57_in = Y57_next;
		Y58_in = Y58_next;
		Y59_in = Y59_next;
		Y60_in = Y60_next;
		Y61_in = Y61_next;
		Y62_in = Y62_next;
		Y63_in = Y63_next;
		Y64_in = Y64_next;
		Y65_in = Y65_next;
		Y66_in = Y66_next;
		Y67_in = Y67_next;
		Y68_in = Y68_next;
		Y69_in = Y69_next;
		Y70_in = Y70_next;
		Y71_in = Y71_next;
		Y72_in = Y72_next;
		Y73_in = Y73_next;
		Y74_in = Y74_next;
		Y75_in = Y75_next;
		Y76_in = Y76_next;
		Y77_in = Y77_next;
		Y78_in = Y78_next;
		Y79_in = Y79_next;
		Y80_in = Y80_next;
		Y81_in = Y81_next;
		Y82_in = Y82_next;
		Y83_in = Y83_next;
		Y84_in = Y84_next;
		Y85_in = Y85_next;
		Y86_in = Y86_next;
		Y87_in = Y87_next;
		Y88_in = Y88_next;
		Y89_in = Y89_next;
		Y90_in = Y90_next;
		Y91_in = Y91_next;
		Y92_in = Y92_next;
		Y93_in = Y93_next;
		Y94_in = Y94_next;
		Y95_in = Y95_next;
		Y96_in = Y96_next;
		Y97_in = Y97_next;
		Y98_in = Y98_next;
		Y99_in = Y99_next;
		Y100_in = Y100_next;
		Y101_in = Y101_next;
		Y102_in = Y102_next;
		Y103_in = Y103_next;
		Y104_in = Y104_next;
		Y105_in = Y105_next;
		Y106_in = Y106_next;
		Y107_in = Y107_next;
		Y108_in = Y108_next;
		Y109_in = Y109_next;
		Y110_in = Y110_next;
		Y111_in = Y111_next;
		Y112_in = Y112_next;
		Y113_in = Y113_next;
		Y114_in = Y114_next;
		Y115_in = Y115_next;
		Y116_in = Y116_next;
		Y117_in = Y117_next;
		Y118_in = Y118_next;
		Y119_in = Y119_next;
		Y120_in = Y120_next;
		Y121_in = Y121_next;
		Y122_in = Y122_next;
		Y123_in = Y123_next;
		Y124_in = Y124_next;
		Y125_in = Y125_next;
		Y126_in = Y126_next;
		Y127_in = Y127_next;
		Y128_in = Y128_next;
		Y129_in = Y129_next;
		Y130_in = Y130_next;
		Y131_in = Y131_next;
		Y132_in = Y132_next;
		Y133_in = Y133_next;
		Y134_in = Y134_next;
		Y135_in = Y135_next;
		Y136_in = Y136_next;
		Y137_in = Y137_next;
		Y138_in = Y138_next;
		Y139_in = Y139_next;
		Y140_in = Y140_next;
		Y141_in = Y141_next;
		Y142_in = Y142_next;
		Y143_in = Y143_next;
		Y144_in = Y144_next;
		Y145_in = Y145_next;
		Y146_in = Y146_next;
		Y147_in = Y147_next;
		Y148_in = Y148_next;
		Y149_in = Y149_next;
		Y150_in = Y150_next;
		Y151_in = Y151_next;
		Y152_in = Y152_next;
		Y153_in = Y153_next;
		Y154_in = Y154_next;
		Y155_in = Y155_next;
		Y156_in = Y156_next;
		Y157_in = Y157_next;
		Y158_in = Y158_next;
		Y159_in = Y159_next;
		Y160_in = Y160_next;
		Y161_in = Y161_next;
		Y162_in = Y162_next;
		Y163_in = Y163_next;
		Y164_in = Y164_next;
		Y165_in = Y165_next;
		Y166_in = Y166_next;
		Y167_in = Y167_next;
		Y168_in = Y168_next;
		Y169_in = Y169_next;
		Y170_in = Y170_next;
		Y171_in = Y171_next;
		Y172_in = Y172_next;
		Y173_in = Y173_next;
		Y174_in = Y174_next;
		Y175_in = Y175_next;
		Y176_in = Y176_next;
		Y177_in = Y177_next;
		Y178_in = Y178_next;
		Y179_in = Y179_next;
		Y180_in = Y180_next;
		Y181_in = Y181_next;
		Y182_in = Y182_next;
		Y183_in = Y183_next;
		Y184_in = Y184_next;
		Y185_in = Y185_next;
		Y186_in = Y186_next;
		Y187_in = Y187_next;
		Y188_in = Y188_next;
		Y189_in = Y189_next;
		Y190_in = Y190_next;
		Y191_in = Y191_next;
		Y192_in = Y192_next;
		Y193_in = Y193_next;
		Y194_in = Y194_next;
		Y195_in = Y195_next;
		Y196_in = Y196_next;
		Y197_in = Y197_next;
		Y198_in = Y198_next;
		Y199_in = Y199_next;
		Y200_in = Y200_next;
		Y201_in = Y201_next;
		Y202_in = Y202_next;
		Y203_in = Y203_next;
		Y204_in = Y204_next;
		Y205_in = Y205_next;
		Y206_in = Y206_next;
		Y207_in = Y207_next;
		Y208_in = Y208_next;
		Y209_in = Y209_next;
		Y210_in = Y210_next;
		Y211_in = Y211_next;
		Y212_in = Y212_next;
		Y213_in = Y213_next;
		Y214_in = Y214_next;
		Y215_in = Y215_next;
		Y216_in = Y216_next;
		Y217_in = Y217_next;
		Y218_in = Y218_next;
		Y219_in = Y219_next;
		Y220_in = Y220_next;
		Y221_in = Y221_next;
		Y222_in = Y222_next;
		Y223_in = Y223_next;
		Y224_in = Y224_next;
		Y225_in = Y225_next;
		Y226_in = Y226_next;
		Y227_in = Y227_next;
		Y228_in = Y228_next;
		Y229_in = Y229_next;
		Y230_in = Y230_next;
		Y231_in = Y231_next;
		Y232_in = Y232_next;
		Y233_in = Y233_next;
		Y234_in = Y234_next;
		Y235_in = Y235_next;
		Y236_in = Y236_next;
		Y237_in = Y237_next;
		Y238_in = Y238_next;
		Y239_in = Y239_next;
		Y240_in = Y240_next;
		Y241_in = Y241_next;
		Y242_in = Y242_next;
		Y243_in = Y243_next;
		Y244_in = Y244_next;
		Y245_in = Y245_next;
		Y246_in = Y246_next;
		Y247_in = Y247_next;
		Y248_in = Y248_next;
		Y249_in = Y249_next;
		Y250_in = Y250_next;
		Y251_in = Y251_next;
		Y252_in = Y252_next;
		Y253_in = Y253_next;
		Y254_in = Y254_next;
		Y255_in = Y255_next;
		Y256_in = Y256_next;		  
	end else begin
		Initial_X = Initial_X_in;
		initial_flag = 1'b0;
	end
	
	U1 <= `WIDTH'b0;
	U2 <= `WIDTH'b0;
	U3 <= `WIDTH'b0;
	U4 <= `WIDTH'b0;
	U5 <= U1_in;
	U6 <= U2_in;
	U7 <= `WIDTH'b0;
	U8 <= U17_in;
	U9 <= U18_in;
  
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y1_in;
    Y6 <= Y2_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y17_in;
    Y9 <= Y18_in;   

    
  end else if (counter == `COUNTER_WIDTH'b01) begin // 2
    
    Y1_next <= onebyoneout;
    
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U1_in;
    U5 <= U2_in;
    U6 <= U3_in;
    U7 <= U17_in;
    U8 <= U18_in;
    U9 <= U19_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y1_in;
    Y5 <= Y2_in;
    Y6 <= Y3_in;
    Y7 <= Y17_in;
    Y8 <= Y18_in;
    Y9 <= Y19_in; 
           

  end else if (counter == `COUNTER_WIDTH'b10) begin // 3
  
    Y2_next <= onebyoneout; 
      
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U2_in;
    U5 <= U3_in;
    U6 <= U4_in;
    U7 <= U18_in;
    U8 <= U19_in;
    U9 <= U20_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y2_in;
    Y5 <= Y3_in;
    Y6 <= Y4_in;
    Y7 <= Y18_in;
    Y8 <= Y19_in;
    Y9 <= Y20_in;
      

  end else if (counter == `COUNTER_WIDTH'b11) begin // 4
  
    Y3_next <= onebyoneout; 
      
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U3_in;
    U5 <= U4_in;
    U6 <= U5_in;
    U7 <= U19_in;
    U8 <= U20_in;
    U9 <= U21_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y3_in;
    Y5 <= Y4_in;
    Y6 <= Y5_in;
    Y7 <= Y19_in;
    Y8 <= Y20_in;
    Y9 <= Y21_in;
       

  end else if (counter == `COUNTER_WIDTH'b100) begin // 5
  
    Y4_next <= onebyoneout;
    
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U4_in;
    U5 <= U5_in;
    U6 <= U6_in;
    U7 <= U20_in;
    U8 <= U21_in;
    U9 <= U22_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y4_in;
    Y5 <= Y5_in;
    Y6 <= Y6_in;
    Y7 <= Y20_in;
    Y8 <= Y21_in;
    Y9 <= Y22_in;
    
    
  end else if (counter == `COUNTER_WIDTH'b101) begin // 6
  
    Y5_next <= onebyoneout;  
  
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U5_in;
    U5 <= U6_in;
    U6 <= U7_in;
    U7 <= U21_in;
    U8 <= U22_in;
    U9 <= U23_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y5_in;
    Y5 <= Y6_in;
    Y6 <= Y7_in;
    Y7 <= Y21_in;
    Y8 <= Y22_in;
    Y9 <= Y23_in;
    

  end else if (counter == `COUNTER_WIDTH'b110) begin // 7
  
    Y6_next <= onebyoneout;
    
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U6_in;
    U5 <= U7_in;
    U6 <= U8_in;
    U7 <= U22_in;
    U8 <= U23_in;
    U9 <= U24_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y6_in;
    Y5 <= Y7_in;
    Y6 <= Y8_in;
    Y7 <= Y22_in;
    Y8 <= Y23_in;
    Y9 <= Y24_in;
    
    
  end else if (counter == `COUNTER_WIDTH'b111) begin // 8

    Y7_next <= onebyoneout;
    
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U7_in;
    U5 <= U8_in;
    U6 <= U9_in;
    U7 <= U23_in;
    U8 <= U24_in;
    U9 <= U25_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y7_in;
    Y5 <= Y8_in;
    Y6 <= Y9_in;
    Y7 <= Y23_in;
    Y8 <= Y24_in;
    Y9 <= Y25_in;
    
    

  end else if (counter == `COUNTER_WIDTH'b1000) begin // 9
 
    Y8_next <= onebyoneout;
     
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U8_in;
    U5 <= U9_in;
    U6 <= U10_in;
    U7 <= U24_in;
    U8 <= U25_in;
    U9 <= U26_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y8_in;
    Y5 <= Y9_in;
    Y6 <= Y10_in;
    Y7 <= Y24_in;
    Y8 <= Y25_in;
    Y9 <= Y26_in;
    
    
 
  end else if (counter == `COUNTER_WIDTH'b1001) begin // 10

    Y9_next <= onebyoneout;
     
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U9_in;
    U5 <= U10_in;
    U6 <= U11_in;
    U7 <= U25_in;
    U8 <= U26_in;
    U9 <= U27_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y9_in;
    Y5 <= Y10_in;
    Y6 <= Y11_in;
    Y7 <= Y25_in;
    Y8 <= Y26_in;
    Y9 <= Y27_in;
    

  end else if (counter == `COUNTER_WIDTH'b1010) begin // 11

    Y10_next <= onebyoneout;
      
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U10_in;
    U5 <= U11_in;
    U6 <= U12_in;
    U7 <= U26_in;
    U8 <= U27_in;
    U9 <= U28_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y10_in;
    Y5 <= Y11_in;
    Y6 <= Y12_in;
    Y7 <= Y26_in;
    Y8 <= Y27_in;
    Y9 <= Y28_in;
    
    

  end else if (counter == `COUNTER_WIDTH'b1011) begin // 12

    Y11_next <= onebyoneout;
      
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U11_in;
    U5 <= U12_in;
    U6 <= U13_in;
    U7 <= U27_in;
    U8 <= U28_in;
    U9 <= U29_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y11_in;
    Y5 <= Y12_in;
    Y6 <= Y13_in;
    Y7 <= Y27_in;
    Y8 <= Y28_in;
    Y9 <= Y29_in;
    

  end else if (counter == `COUNTER_WIDTH'b1100) begin // 13

    Y12_next <= onebyoneout;
      
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U12_in;
    U5 <= U13_in;
    U6 <= U14_in;
    U7 <= U28_in;
    U8 <= U29_in;
    U9 <= U30_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y12_in;
    Y5 <= Y13_in;
    Y6 <= Y14_in;
    Y7 <= Y28_in;
    Y8 <= Y29_in;
    Y9 <= Y30_in;
    

  end else if (counter == `COUNTER_WIDTH'b1101) begin // 14

    Y13_next <= onebyoneout;
      
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U13_in;
    U5 <= U14_in;
    U6 <= U15_in;
    U7 <= U29_in;
    U8 <= U30_in;
    U9 <= U31_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y13_in;
    Y5 <= Y14_in;
    Y6 <= Y15_in;
    Y7 <= Y29_in;
    Y8 <= Y30_in;
    Y9 <= Y31_in;
    
    

  end else if (counter == `COUNTER_WIDTH'b1110) begin // 15
 
    Y14_next <= onebyoneout;
      
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U14_in;
    U5 <= U15_in;
    U6 <= U16_in;
    U7 <= U30_in;
    U8 <= U31_in;
    U9 <= U32_in;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y14_in;
    Y5 <= Y15_in;
    Y6 <= Y16_in;
    Y7 <= Y30_in;
    Y8 <= Y31_in;
    Y9 <= Y32_in;
    

  end else if (counter == `COUNTER_WIDTH'b1111) begin // 16
  
    Y15_next <= onebyoneout;
    
    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U15_in;
    U5 <= U16_in;
    U6 <= `WIDTH'b0;
    U7 <= U31_in;
    U8 <= U32_in;
    U9 <= `WIDTH'b0;
    
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y15_in;
    Y5 <= Y16_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y31_in;
    Y8 <= Y32_in;
    Y9 <= {(2 * `WIDTH){1'b0}}; 
      
// 5 bits    
  end else if (counter == `COUNTER_WIDTH'b10000) begin // 17
  
    Y16_next <= onebyoneout;
  
    U1 <= `WIDTH'b0;
	U2 <= U1_in;
	U3 <= U2_in;
	U4 <= `WIDTH'b0;
	U5 <= U17_in;
	U6 <= U18_in;
	U7 <= `WIDTH'b0;
	U8 <= U33_in;
	U9 <= U34_in;
  
    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y1_in;
    Y3 <= Y2_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y17_in;
    Y6 <= Y18_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y33_in;
    Y9 <= Y34_in; 
    
  end else if (counter == `COUNTER_WIDTH'b10001) begin // 18
  
    Y17_next <= onebyoneout;

    U1 <= U1_in;
    U2 <= U2_in;
    U3 <= U3_in;
    U4 <= U17_in;
    U5 <= U18_in;
    U6 <= U19_in;
    U7 <= U33_in;
    U8 <= U34_in;
    U9 <= U35_in;


    Y1 <= Y1_in;
    Y2 <= Y2_in;
    Y3 <= Y3_in;
    Y4 <= Y17_in;
    Y5 <= Y18_in;
    Y6 <= Y19_in;
    Y7 <= Y33_in;
    Y8 <= Y34_in;
    Y9 <= Y35_in;
    
  end else if (counter == `COUNTER_WIDTH'b10010) begin // 19
    
    Y18_next <= onebyoneout;
  
	U1 <= U2_in;
	U2 <= U3_in;
	U3 <= U4_in;
	U4 <= U18_in;
	U5 <= U19_in;
	U6 <= U20_in;
	U7 <= U34_in;
	U8 <= U35_in;
	U9 <= U36_in;
  
    Y1 <= Y2_in;
    Y2 <= Y3_in;
    Y3 <= Y4_in;
    Y4 <= Y18_in;
    Y5 <= Y19_in;
    Y6 <= Y20_in;
    Y7 <= Y34_in;
    Y8 <= Y35_in;
    Y9 <= Y36_in;
    
  end else if (counter == `COUNTER_WIDTH'b10011) begin // 20
      
    Y19_next <= onebyoneout;
  
    U1 <= U3_in;
	U2 <= U4_in;
	U3 <= U5_in;
	U4 <= U19_in;
	U5 <= U20_in;
	U6 <= U21_in;
	U7 <= U35_in;
	U8 <= U36_in;
	U9 <= U37_in;
  
    Y1 <= Y3_in;
    Y2 <= Y4_in;
    Y3 <= Y5_in;
    Y4 <= Y19_in;
    Y5 <= Y20_in;
    Y6 <= Y21_in;
    Y7 <= Y35_in;
    Y8 <= Y36_in;
    Y9 <= Y37_in;
 
  end else if (counter == `COUNTER_WIDTH'b10100) begin // 21
        
    Y20_next <= onebyoneout;
  
    U1 <= U4_in;
	U2 <= U5_in;
	U3 <= U6_in;
	U4 <= U20_in;
	U5 <= U21_in;
	U6 <= U22_in;
	U7 <= U36_in;
	U8 <= U37_in;
	U9 <= U38_in;
  
    Y1 <= Y4_in;
    Y2 <= Y5_in;
    Y3 <= Y6_in;
    Y4 <= Y20_in;
    Y5 <= Y21_in;
    Y6 <= Y22_in;
    Y7 <= Y36_in;
    Y8 <= Y37_in;
    Y9 <= Y38_in;
 
  end else if (counter == `COUNTER_WIDTH'b10101) begin // 22
          
    Y21_next <= onebyoneout;
  
    U1 <= U5_in;
	U2 <= U6_in;
	U3 <= U7_in;
	U4 <= U21_in;
	U5 <= U22_in;
	U6 <= U23_in;
	U7 <= U37_in;
	U8 <= U38_in;
	U9 <= U39_in;
  
    Y1 <= Y5_in;
    Y2 <= Y6_in;
    Y3 <= Y7_in;
    Y4 <= Y21_in;
    Y5 <= Y22_in;
    Y6 <= Y23_in;
    Y7 <= Y37_in;
    Y8 <= Y38_in;
    Y9 <= Y39_in;
 
  end else if (counter == `COUNTER_WIDTH'b10110) begin // 23
 
    Y22_next <= onebyoneout;

    U1 <= U6_in;
    U2 <= U7_in;
    U3 <= U8_in;
    U4 <= U22_in;
    U5 <= U23_in;
    U6 <= U24_in;
    U7 <= U38_in;
    U8 <= U39_in;
    U9 <= U40_in;
    
    Y1 <= Y6_in;
    Y2 <= Y7_in;
    Y3 <= Y8_in;
    Y4 <= Y22_in;
    Y5 <= Y23_in;
    Y6 <= Y24_in;
    Y7 <= Y38_in;
    Y8 <= Y39_in;
    Y9 <= Y40_in;

  end else if (counter == `COUNTER_WIDTH'b10111) begin // 24

    Y23_next <= onebyoneout;

    U1 <= U7_in;
    U2 <= U8_in;
    U3 <= U9_in;
    U4 <= U23_in;
    U5 <= U24_in;
    U6 <= U25_in;
    U7 <= U39_in;
    U8 <= U40_in;
    U9 <= U41_in;

    Y1 <= Y7_in;
    Y2 <= Y8_in;
    Y3 <= Y9_in;
    Y4 <= Y23_in;
    Y5 <= Y24_in;
    Y6 <= Y25_in;
    Y7 <= Y39_in;
    Y8 <= Y40_in;
    Y9 <= Y41_in;
  
  end else if (counter == `COUNTER_WIDTH'b11000) begin // 25
  
    Y24_next <= onebyoneout;

    U1 <= U8_in;
    U2 <= U9_in;
    U3 <= U10_in;
    U4 <= U24_in;
    U5 <= U25_in;
    U6 <= U26_in;
    U7 <= U40_in;
    U8 <= U41_in;
    U9 <= U42_in;

    Y1 <= Y8_in;
    Y2 <= Y9_in;
    Y3 <= Y10_in;
    Y4 <= Y24_in;
    Y5 <= Y25_in;
    Y6 <= Y26_in;
    Y7 <= Y40_in;
    Y8 <= Y41_in;
    Y9 <= Y42_in;

  end else if (counter == `COUNTER_WIDTH'b11001) begin // 26
  
  	Y25_next <= onebyoneout;

    U1 <= U9_in;
    U2 <= U10_in;
    U3 <= U11_in;
    U4 <= U25_in;
    U5 <= U26_in;
    U6 <= U27_in;
    U7 <= U41_in;
    U8 <= U42_in;
    U9 <= U43_in;

    Y1 <= Y9_in;
    Y2 <= Y10_in;
    Y3 <= Y11_in;
    Y4 <= Y25_in;
    Y5 <= Y26_in;
    Y6 <= Y27_in;
    Y7 <= Y41_in;
    Y8 <= Y42_in;
    Y9 <= Y43_in;

  end else if (counter == `COUNTER_WIDTH'b11010) begin // 27
  
    Y26_next <= onebyoneout;

    U1 <= U10_in;
    U2 <= U11_in;
    U3 <= U12_in;
    U4 <= U26_in;
    U5 <= U27_in;
    U6 <= U28_in;
    U7 <= U42_in;
    U8 <= U43_in;
    U9 <= U44_in;


    Y1 <= Y10_in;
    Y2 <= Y11_in;
    Y3 <= Y12_in;
    Y4 <= Y26_in;
    Y5 <= Y27_in;
    Y6 <= Y28_in;
    Y7 <= Y42_in;
    Y8 <= Y43_in;
    Y9 <= Y44_in;

  end else if (counter == `COUNTER_WIDTH'b11011) begin // 28
  
    Y27_next <= onebyoneout;

    U1 <= U11_in;
    U2 <= U12_in;
    U3 <= U13_in;
    U4 <= U27_in;
    U5 <= U28_in;
    U6 <= U29_in;
    U7 <= U43_in;
    U8 <= U44_in;
    U9 <= U45_in;

    Y1 <= Y11_in;
    Y2 <= Y12_in;
    Y3 <= Y13_in;
    Y4 <= Y27_in;
    Y5 <= Y28_in;
    Y6 <= Y29_in;
    Y7 <= Y43_in;
    Y8 <= Y44_in;
    Y9 <= Y45_in;

  end else if (counter == `COUNTER_WIDTH'b11100) begin // 29
  
    Y28_next <= onebyoneout;

    U1 <= U12_in;
    U2 <= U13_in;
    U3 <= U14_in;
    U4 <= U28_in;
    U5 <= U29_in;
    U6 <= U30_in;
    U7 <= U44_in;
    U8 <= U45_in;
    U9 <= U46_in;

    Y1 <= Y12_in;
    Y2 <= Y13_in;
    Y3 <= Y14_in;
    Y4 <= Y28_in;
    Y5 <= Y29_in;
    Y6 <= Y30_in;
    Y7 <= Y44_in;
    Y8 <= Y45_in;
    Y9 <= Y46_in;


  end else if (counter == `COUNTER_WIDTH'b11101) begin // 30
  
    Y29_next <= onebyoneout;

    U1 <= U13_in;
    U2 <= U14_in;
    U3 <= U15_in;
    U4 <= U29_in;
    U5 <= U30_in;
    U6 <= U31_in;
    U7 <= U45_in;
    U8 <= U46_in;
    U9 <= U47_in;


    Y1 <= Y13_in;
    Y2 <= Y14_in;
    Y3 <= Y15_in;
    Y4 <= Y29_in;
    Y5 <= Y30_in;
    Y6 <= Y31_in;
    Y7 <= Y45_in;
    Y8 <= Y46_in;
    Y9 <= Y47_in;

  end else if (counter == `COUNTER_WIDTH'b11110) begin // 31
  
    Y30_next <= onebyoneout;

    U1 <= U14_in;
    U2 <= U15_in;
    U3 <= U16_in;
    U4 <= U30_in;
    U5 <= U31_in;
    U6 <= U32_in;
    U7 <= U46_in;
    U8 <= U47_in;
    U9 <= U48_in;


    Y1 <= Y14_in;
    Y2 <= Y15_in;
    Y3 <= Y16_in;
    Y4 <= Y30_in;
    Y5 <= Y31_in;
    Y6 <= Y32_in;
    Y7 <= Y46_in;
    Y8 <= Y47_in;
    Y9 <= Y48_in;

  end else if (counter == `COUNTER_WIDTH'b11111) begin // 32
  
    Y31_next <= onebyoneout;
    
    U1 <= U15_in;
    U2 <= U16_in;
    U3 <= `WIDTH'b0;
    U4 <= U31_in;
    U5 <= U32_in;
    U6 <= `WIDTH'b0;
    U7 <= U47_in;
    U8 <= U48_in;
    U9 <= `WIDTH'b0;
    
    Y1 <= Y15_in;
    Y2 <= Y16_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y31_in;
    Y5 <= Y32_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y47_in;
    Y8 <= Y48_in;
    Y9 <= {(2 * `WIDTH){1'b0}}; 
      
// 6 bits
  end else if (counter == `COUNTER_WIDTH'b100000) begin
  end else if (counter == `COUNTER_WIDTH'b100001) begin
  end else if (counter == `COUNTER_WIDTH'b100010) begin
  end else if (counter == `COUNTER_WIDTH'b100011) begin
  end else if (counter == `COUNTER_WIDTH'b100100) begin
  end else if (counter == `COUNTER_WIDTH'b100101) begin
  end else if (counter == `COUNTER_WIDTH'b100110) begin
  end else if (counter == `COUNTER_WIDTH'b100111) begin
  end else if (counter == `COUNTER_WIDTH'b101000) begin
  end else if (counter == `COUNTER_WIDTH'b101001) begin
  end else if (counter == `COUNTER_WIDTH'b101010) begin
  end else if (counter == `COUNTER_WIDTH'b101011) begin
  end else if (counter == `COUNTER_WIDTH'b101100) begin
  end else if (counter == `COUNTER_WIDTH'b101101) begin
  end else if (counter == `COUNTER_WIDTH'b101110) begin
  end else if (counter == `COUNTER_WIDTH'b101111) begin

  end else if (counter == `COUNTER_WIDTH'b110000) begin
  end else if (counter == `COUNTER_WIDTH'b110001) begin
  end else if (counter == `COUNTER_WIDTH'b110010) begin
  end else if (counter == `COUNTER_WIDTH'b110011) begin
  end else if (counter == `COUNTER_WIDTH'b110100) begin
  end else if (counter == `COUNTER_WIDTH'b110101) begin
  end else if (counter == `COUNTER_WIDTH'b110110) begin
  end else if (counter == `COUNTER_WIDTH'b110111) begin
  end else if (counter == `COUNTER_WIDTH'b111000) begin
  end else if (counter == `COUNTER_WIDTH'b111001) begin
  end else if (counter == `COUNTER_WIDTH'b111010) begin
  end else if (counter == `COUNTER_WIDTH'b111011) begin
  end else if (counter == `COUNTER_WIDTH'b111100) begin
  end else if (counter == `COUNTER_WIDTH'b111101) begin
  end else if (counter == `COUNTER_WIDTH'b111110) begin
  end else if (counter == `COUNTER_WIDTH'b111111) begin
// 7 bits
  end else if (counter == `COUNTER_WIDTH'b1000000) begin
  end else if (counter == `COUNTER_WIDTH'b1000001) begin
  end else if (counter == `COUNTER_WIDTH'b1000010) begin
  end else if (counter == `COUNTER_WIDTH'b1000011) begin
  end else if (counter == `COUNTER_WIDTH'b1000100) begin
  end else if (counter == `COUNTER_WIDTH'b1000101) begin
  end else if (counter == `COUNTER_WIDTH'b1000110) begin
  end else if (counter == `COUNTER_WIDTH'b1000111) begin
  end else if (counter == `COUNTER_WIDTH'b1001000) begin
  end else if (counter == `COUNTER_WIDTH'b1001001) begin
  end else if (counter == `COUNTER_WIDTH'b1001010) begin
  end else if (counter == `COUNTER_WIDTH'b1001011) begin
  end else if (counter == `COUNTER_WIDTH'b1001100) begin
  end else if (counter == `COUNTER_WIDTH'b1001101) begin
  end else if (counter == `COUNTER_WIDTH'b1001110) begin
  end else if (counter == `COUNTER_WIDTH'b1001111) begin

  end else if (counter == `COUNTER_WIDTH'b1010000) begin
  end else if (counter == `COUNTER_WIDTH'b1010001) begin
  end else if (counter == `COUNTER_WIDTH'b1010010) begin
  end else if (counter == `COUNTER_WIDTH'b1010011) begin
  end else if (counter == `COUNTER_WIDTH'b1010100) begin
  end else if (counter == `COUNTER_WIDTH'b1010101) begin
  end else if (counter == `COUNTER_WIDTH'b1010110) begin
  end else if (counter == `COUNTER_WIDTH'b1010111) begin
  end else if (counter == `COUNTER_WIDTH'b1011000) begin
  end else if (counter == `COUNTER_WIDTH'b1011001) begin
  end else if (counter == `COUNTER_WIDTH'b1011010) begin
  end else if (counter == `COUNTER_WIDTH'b1011011) begin
  end else if (counter == `COUNTER_WIDTH'b1011100) begin
  end else if (counter == `COUNTER_WIDTH'b1011101) begin
  end else if (counter == `COUNTER_WIDTH'b1011110) begin
  end else if (counter == `COUNTER_WIDTH'b1011111) begin

  end else if (counter == `COUNTER_WIDTH'b1100000) begin
  end else if (counter == `COUNTER_WIDTH'b1100001) begin
  end else if (counter == `COUNTER_WIDTH'b1100010) begin
  end else if (counter == `COUNTER_WIDTH'b1100011) begin
  end else if (counter == `COUNTER_WIDTH'b1100100) begin
  end else if (counter == `COUNTER_WIDTH'b1100101) begin
  end else if (counter == `COUNTER_WIDTH'b1100110) begin
  end else if (counter == `COUNTER_WIDTH'b1100111) begin
  end else if (counter == `COUNTER_WIDTH'b1101000) begin
  end else if (counter == `COUNTER_WIDTH'b1101001) begin
  end else if (counter == `COUNTER_WIDTH'b1101010) begin
  end else if (counter == `COUNTER_WIDTH'b1101011) begin
  end else if (counter == `COUNTER_WIDTH'b1101100) begin
  end else if (counter == `COUNTER_WIDTH'b1101101) begin
  end else if (counter == `COUNTER_WIDTH'b1101110) begin
  end else if (counter == `COUNTER_WIDTH'b1101111) begin

  end else if (counter == `COUNTER_WIDTH'b1110000) begin
  end else if (counter == `COUNTER_WIDTH'b1110001) begin
  end else if (counter == `COUNTER_WIDTH'b1110010) begin
  end else if (counter == `COUNTER_WIDTH'b1110011) begin
  end else if (counter == `COUNTER_WIDTH'b1110100) begin
  end else if (counter == `COUNTER_WIDTH'b1110101) begin
  end else if (counter == `COUNTER_WIDTH'b1110110) begin
  end else if (counter == `COUNTER_WIDTH'b1110111) begin
  end else if (counter == `COUNTER_WIDTH'b1111000) begin
  end else if (counter == `COUNTER_WIDTH'b1111001) begin
  end else if (counter == `COUNTER_WIDTH'b1111010) begin
  end else if (counter == `COUNTER_WIDTH'b1111011) begin
  end else if (counter == `COUNTER_WIDTH'b1111100) begin
  end else if (counter == `COUNTER_WIDTH'b1111101) begin
  end else if (counter == `COUNTER_WIDTH'b1111110) begin
  end else if (counter == `COUNTER_WIDTH'b1111111) begin
// 8 bits
  end else if (counter == `COUNTER_WIDTH'b10000000) begin
  end else if (counter == `COUNTER_WIDTH'b10000001) begin
  end else if (counter == `COUNTER_WIDTH'b10000010) begin
  end else if (counter == `COUNTER_WIDTH'b10000011) begin
  end else if (counter == `COUNTER_WIDTH'b10000100) begin
  end else if (counter == `COUNTER_WIDTH'b10000101) begin
  end else if (counter == `COUNTER_WIDTH'b10000110) begin
  end else if (counter == `COUNTER_WIDTH'b10000111) begin
  end else if (counter == `COUNTER_WIDTH'b10001000) begin
  end else if (counter == `COUNTER_WIDTH'b10001001) begin
  end else if (counter == `COUNTER_WIDTH'b10001010) begin
  end else if (counter == `COUNTER_WIDTH'b10001011) begin
  end else if (counter == `COUNTER_WIDTH'b10001100) begin
  end else if (counter == `COUNTER_WIDTH'b10001101) begin
  end else if (counter == `COUNTER_WIDTH'b10001110) begin
  end else if (counter == `COUNTER_WIDTH'b10001111) begin

  end else if (counter == `COUNTER_WIDTH'b10010000) begin
  end else if (counter == `COUNTER_WIDTH'b10010001) begin
  end else if (counter == `COUNTER_WIDTH'b10010010) begin
  end else if (counter == `COUNTER_WIDTH'b10010011) begin
  end else if (counter == `COUNTER_WIDTH'b10010100) begin
  end else if (counter == `COUNTER_WIDTH'b10010101) begin
  end else if (counter == `COUNTER_WIDTH'b10010110) begin
  end else if (counter == `COUNTER_WIDTH'b10010111) begin
  end else if (counter == `COUNTER_WIDTH'b10011000) begin
  end else if (counter == `COUNTER_WIDTH'b10011001) begin
  end else if (counter == `COUNTER_WIDTH'b10011010) begin
  end else if (counter == `COUNTER_WIDTH'b10011011) begin
  end else if (counter == `COUNTER_WIDTH'b10011100) begin
  end else if (counter == `COUNTER_WIDTH'b10011101) begin
  end else if (counter == `COUNTER_WIDTH'b10011110) begin
  end else if (counter == `COUNTER_WIDTH'b10011111) begin

  end else if (counter == `COUNTER_WIDTH'b10100000) begin
  end else if (counter == `COUNTER_WIDTH'b10100001) begin
  end else if (counter == `COUNTER_WIDTH'b10100010) begin
  end else if (counter == `COUNTER_WIDTH'b10100011) begin
  end else if (counter == `COUNTER_WIDTH'b10100100) begin
  end else if (counter == `COUNTER_WIDTH'b10100101) begin
  end else if (counter == `COUNTER_WIDTH'b10100110) begin
  end else if (counter == `COUNTER_WIDTH'b10100111) begin
  end else if (counter == `COUNTER_WIDTH'b10101000) begin
  end else if (counter == `COUNTER_WIDTH'b10101001) begin
  end else if (counter == `COUNTER_WIDTH'b10101010) begin
  end else if (counter == `COUNTER_WIDTH'b10101011) begin
  end else if (counter == `COUNTER_WIDTH'b10101100) begin
  end else if (counter == `COUNTER_WIDTH'b10101101) begin
  end else if (counter == `COUNTER_WIDTH'b10101110) begin
  end else if (counter == `COUNTER_WIDTH'b10101111) begin

  end else if (counter == `COUNTER_WIDTH'b10110000) begin
  end else if (counter == `COUNTER_WIDTH'b10110001) begin
  end else if (counter == `COUNTER_WIDTH'b10110010) begin
  end else if (counter == `COUNTER_WIDTH'b10110011) begin
  end else if (counter == `COUNTER_WIDTH'b10110100) begin
  end else if (counter == `COUNTER_WIDTH'b10110101) begin
  end else if (counter == `COUNTER_WIDTH'b10110110) begin
  end else if (counter == `COUNTER_WIDTH'b10110111) begin
  end else if (counter == `COUNTER_WIDTH'b10111000) begin
  end else if (counter == `COUNTER_WIDTH'b10111001) begin
  end else if (counter == `COUNTER_WIDTH'b10111010) begin
  end else if (counter == `COUNTER_WIDTH'b10111011) begin
  end else if (counter == `COUNTER_WIDTH'b10111100) begin
  end else if (counter == `COUNTER_WIDTH'b10111101) begin
  end else if (counter == `COUNTER_WIDTH'b10111110) begin
  end else if (counter == `COUNTER_WIDTH'b10111111) begin

  end else if (counter == `COUNTER_WIDTH'b11000000) begin
  end else if (counter == `COUNTER_WIDTH'b11000001) begin
  end else if (counter == `COUNTER_WIDTH'b11000010) begin
  end else if (counter == `COUNTER_WIDTH'b11000011) begin
  end else if (counter == `COUNTER_WIDTH'b11000100) begin
  end else if (counter == `COUNTER_WIDTH'b11000101) begin
  end else if (counter == `COUNTER_WIDTH'b11000110) begin
  end else if (counter == `COUNTER_WIDTH'b11000111) begin
  end else if (counter == `COUNTER_WIDTH'b11001000) begin
  end else if (counter == `COUNTER_WIDTH'b11001001) begin
  end else if (counter == `COUNTER_WIDTH'b11001010) begin
  end else if (counter == `COUNTER_WIDTH'b11001011) begin
  end else if (counter == `COUNTER_WIDTH'b11001100) begin
  end else if (counter == `COUNTER_WIDTH'b11001101) begin
  end else if (counter == `COUNTER_WIDTH'b11001110) begin
  end else if (counter == `COUNTER_WIDTH'b11001111) begin

  end else if (counter == `COUNTER_WIDTH'b11010000) begin
  end else if (counter == `COUNTER_WIDTH'b11010001) begin
  end else if (counter == `COUNTER_WIDTH'b11010010) begin
  end else if (counter == `COUNTER_WIDTH'b11010011) begin
  end else if (counter == `COUNTER_WIDTH'b11010100) begin
  end else if (counter == `COUNTER_WIDTH'b11010101) begin
  end else if (counter == `COUNTER_WIDTH'b11010110) begin
  end else if (counter == `COUNTER_WIDTH'b11010111) begin
  end else if (counter == `COUNTER_WIDTH'b11011000) begin
  end else if (counter == `COUNTER_WIDTH'b11011001) begin
  end else if (counter == `COUNTER_WIDTH'b11011010) begin
  end else if (counter == `COUNTER_WIDTH'b11011011) begin
  end else if (counter == `COUNTER_WIDTH'b11011100) begin
  end else if (counter == `COUNTER_WIDTH'b11011101) begin
  end else if (counter == `COUNTER_WIDTH'b11011110) begin
  end else if (counter == `COUNTER_WIDTH'b11011111) begin

  end else if (counter == `COUNTER_WIDTH'b11100000) begin
  end else if (counter == `COUNTER_WIDTH'b11100001) begin
  end else if (counter == `COUNTER_WIDTH'b11100010) begin
  end else if (counter == `COUNTER_WIDTH'b11100011) begin
  end else if (counter == `COUNTER_WIDTH'b11100100) begin
  end else if (counter == `COUNTER_WIDTH'b11100101) begin
  end else if (counter == `COUNTER_WIDTH'b11100110) begin
  end else if (counter == `COUNTER_WIDTH'b11100111) begin
  end else if (counter == `COUNTER_WIDTH'b11101000) begin
  end else if (counter == `COUNTER_WIDTH'b11101001) begin
  end else if (counter == `COUNTER_WIDTH'b11101010) begin
  end else if (counter == `COUNTER_WIDTH'b11101011) begin
  end else if (counter == `COUNTER_WIDTH'b11101100) begin
  end else if (counter == `COUNTER_WIDTH'b11101101) begin
  end else if (counter == `COUNTER_WIDTH'b11101110) begin
  end else if (counter == `COUNTER_WIDTH'b11101111) begin

  end else if (counter == `COUNTER_WIDTH'b11110000) begin
  end else if (counter == `COUNTER_WIDTH'b11110001) begin
  end else if (counter == `COUNTER_WIDTH'b11110010) begin
  end else if (counter == `COUNTER_WIDTH'b11110011) begin
  end else if (counter == `COUNTER_WIDTH'b11110100) begin
  end else if (counter == `COUNTER_WIDTH'b11110101) begin
  end else if (counter == `COUNTER_WIDTH'b11110110) begin
  end else if (counter == `COUNTER_WIDTH'b11110111) begin
  end else if (counter == `COUNTER_WIDTH'b11111000) begin
  end else if (counter == `COUNTER_WIDTH'b11111001) begin
  end else if (counter == `COUNTER_WIDTH'b11111010) begin
  end else if (counter == `COUNTER_WIDTH'b11111011) begin
  end else if (counter == `COUNTER_WIDTH'b11111100) begin
  end else if (counter == `COUNTER_WIDTH'b11111101) begin
  end else if (counter == `COUNTER_WIDTH'b11111110) begin
  end else if (counter == `COUNTER_WIDTH'b11111111) begin // 256
    
    Y255_next <= onebyoneout;
      
    U1 <= U239_in;
    U2 <= U240_in;
    U3 <= `WIDTH'b0;
    U4 <= U255_in;
    U5 <= U256_in;
    U6 <= `WIDTH'b0;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    Y1 <= Y239_in;
    Y2 <= Y240_in;
    Y3 <= `WIDTH'b0;
    Y4 <= Y255_in;
    Y5 <= Y256_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};
    end
  counter = counter + `COUNTER_WIDTH'b1;
end




onebyone u1(
.A1(A1[`WIDTH - 1:0]),
.A2(A2[`WIDTH - 1:0]),
.A3(A3[`WIDTH - 1:0]),
.A4(A4[`WIDTH - 1:0]),
.A5(A5[`WIDTH - 1:0]),
.A6(A6[`WIDTH - 1:0]),
.A7(A7[`WIDTH - 1:0]),
.A8(A8[`WIDTH - 1:0]),
.A9(A9[`WIDTH - 1:0]),

.B1(B1[`WIDTH - 1:0]),
.B2(B2[`WIDTH - 1:0]),
.B3(B3[`WIDTH - 1:0]),
.B4(B4[`WIDTH - 1:0]),
.B5(B5[`WIDTH - 1:0]),
.B6(B6[`WIDTH - 1:0]),
.B7(B7[`WIDTH - 1:0]),
.B8(B8[`WIDTH - 1:0]),
.B9(B9[`WIDTH - 1:0]),

.U1(U1[`WIDTH - 1:0]),
.U2(U2[`WIDTH - 1:0]),
.U3(U3[`WIDTH - 1:0]),
.U4(U4[`WIDTH - 1:0]),
.U5(U5[`WIDTH - 1:0]),
.U6(U6[`WIDTH - 1:0]),
.U7(U7[`WIDTH - 1:0]),
.U8(U8[`WIDTH - 1:0]),
.U9(U9[`WIDTH - 1:0]),

.Y1(Y1[2 * `WIDTH - 1:0]),
.Y2(Y2[2 * `WIDTH - 1:0]),
.Y3(Y3[2 * `WIDTH - 1:0]),
.Y4(Y4[2 * `WIDTH - 1:0]),
.Y5(Y5[2 * `WIDTH - 1:0]),
.Y6(Y6[2 * `WIDTH - 1:0]),
.Y7(Y7[2 * `WIDTH - 1:0]),
.Y8(Y8[2 * `WIDTH - 1:0]),
.Y9(Y9[2 * `WIDTH - 1:0]),

.I(I[`WIDTH - 1:0]),

.Initial_X(Initial_X[2 * `WIDTH - 1:0]),

.out(onebyoneout[2 * `WIDTH - 1:0])

);

endmodule
