`define WIDTH 9
module CNNsixteenbysixteen (
clk,

Y1_out, Y2_out, Y3_out, Y4_out, Y5_out, Y6_out, Y7_out, Y8_out, Y9_out, Y10_out, Y11_out, Y12_out, Y13_out, Y14_out, Y15_out, Y16_out
  );
	input wire clk;
	wire signed [`WIDTH - 1:0] A1, A2, A3, A4, A5, A6, A7, A8, A9;
	wire signed [`WIDTH - 1:0] B1, B2, B3, B4, B5, B6, B7, B8, B9;
	wire signed [`WIDTH - 1:0] I;
	wire signed [`WIDTH - 1:0] U1_in, U2_in, U3_in, U4_in, U5_in, U6_in, U7_in, U8_in, U9_in, U10_in, U11_in, U12_in, U13_in, U14_in, U15_in, U16_in;
	wire signed [`WIDTH - 1:0] U8_in, U9_in, U10_in, U11_in, U12_in, U13_in, U14_in, U15_in, U16_in, U17_in, U18_in, U19_in, U20_in, U21_in, U22_in, U23_in;
	wire signed [`WIDTH - 1:0] U15_in, U16_in, U17_in, U18_in, U19_in, U20_in, U21_in, U22_in, U23_in, U24_in, U25_in, U26_in, U27_in, U28_in, U29_in, U30_in;
	wire signed [`WIDTH - 1:0] U22_in, U23_in, U24_in, U25_in, U26_in, U27_in, U28_in, U29_in, U30_in, U31_in, U32_in, U33_in, U34_in, U35_in, U36_in, U37_in;
	wire signed [`WIDTH - 1:0] U29_in, U30_in, U31_in, U32_in, U33_in, U34_in, U35_in, U36_in, U37_in, U38_in, U39_in, U40_in, U41_in, U42_in, U43_in, U44_in;
	wire signed [`WIDTH - 1:0] U36_in, U37_in, U38_in, U39_in, U40_in, U41_in, U42_in, U43_in, U44_in, U45_in, U46_in, U47_in, U48_in, U49_in, U50_in, U51_in;
	wire signed [`WIDTH - 1:0] U43_in, U44_in, U45_in, U46_in, U47_in, U48_in, U49_in, U50_in, U51_in, U52_in, U53_in, U54_in, U55_in, U56_in, U57_in, U58_in;
	wire signed [`WIDTH - 1:0] U50_in, U51_in, U52_in, U53_in, U54_in, U55_in, U56_in, U57_in, U58_in, U59_in, U60_in, U61_in, U62_in, U63_in, U64_in, U65_in;
	wire signed [`WIDTH - 1:0] U57_in, U58_in, U59_in, U60_in, U61_in, U62_in, U63_in, U64_in, U65_in, U66_in, U67_in, U68_in, U69_in, U70_in, U71_in, U72_in;
	wire signed [`WIDTH - 1:0] U64_in, U65_in, U66_in, U67_in, U68_in, U69_in, U70_in, U71_in, U72_in, U73_in, U74_in, U75_in, U76_in, U77_in, U78_in, U79_in;
	wire signed [`WIDTH - 1:0] U71_in, U72_in, U73_in, U74_in, U75_in, U76_in, U77_in, U78_in, U79_in, U80_in, U81_in, U82_in, U83_in, U84_in, U85_in, U86_in;
	wire signed [`WIDTH - 1:0] U78_in, U79_in, U80_in, U81_in, U82_in, U83_in, U84_in, U85_in, U86_in, U87_in, U88_in, U89_in, U90_in, U91_in, U92_in, U93_in;
	wire signed [`WIDTH - 1:0] U85_in, U86_in, U87_in, U88_in, U89_in, U90_in, U91_in, U92_in, U93_in, U94_in, U95_in, U96_in, U97_in, U98_in, U99_in, U100_in;
	wire signed [`WIDTH - 1:0] U92_in, U93_in, U94_in, U95_in, U96_in, U97_in, U98_in, U99_in, U100_in, U101_in, U102_in, U103_in, U104_in, U105_in, U106_in, U107_in;
	wire signed [`WIDTH - 1:0] U99_in, U100_in, U101_in, U102_in, U103_in, U104_in, U105_in, U106_in, U107_in, U108_in, U109_in, U110_in, U111_in, U112_in, U113_in, U114_in;
	wire signed [`WIDTH - 1:0] U106_in, U107_in, U108_in, U109_in, U110_in, U111_in, U112_in, U113_in, U114_in, U115_in, U116_in, U117_in, U118_in, U119_in, U120_in, U121_in;
	wire signed [`WIDTH - 1:0] U113_in, U114_in, U115_in, U116_in, U117_in, U118_in, U119_in, U120_in, U121_in, U122_in, U123_in, U124_in, U125_in, U126_in, U127_in, U128_in;
	wire signed [`WIDTH - 1:0] U120_in, U121_in, U122_in, U123_in, U124_in, U125_in, U126_in, U127_in, U128_in, U129_in, U130_in, U131_in, U132_in, U133_in, U134_in, U135_in;
	wire signed [`WIDTH - 1:0] U127_in, U128_in, U129_in, U130_in, U131_in, U132_in, U133_in, U134_in, U135_in, U136_in, U137_in, U138_in, U139_in, U140_in, U141_in, U142_in;
	wire signed [`WIDTH - 1:0] U134_in, U135_in, U136_in, U137_in, U138_in, U139_in, U140_in, U141_in, U142_in, U143_in, U144_in, U145_in, U146_in, U147_in, U148_in, U149_in;
	wire signed [`WIDTH - 1:0] U141_in, U142_in, U143_in, U144_in, U145_in, U146_in, U147_in, U148_in, U149_in, U150_in, U151_in, U152_in, U153_in, U154_in, U155_in, U156_in;
	wire signed [`WIDTH - 1:0] U148_in, U149_in, U150_in, U151_in, U152_in, U153_in, U154_in, U155_in, U156_in, U157_in, U158_in, U159_in, U160_in, U161_in, U162_in, U163_in;
	wire signed [`WIDTH - 1:0] U155_in, U156_in, U157_in, U158_in, U159_in, U160_in, U161_in, U162_in, U163_in, U164_in, U165_in, U166_in, U167_in, U168_in, U169_in, U170_in;
	wire signed [`WIDTH - 1:0] U162_in, U163_in, U164_in, U165_in, U166_in, U167_in, U168_in, U169_in, U170_in, U171_in, U172_in, U173_in, U174_in, U175_in, U176_in, U177_in;
	wire signed [`WIDTH - 1:0] U169_in, U170_in, U171_in, U172_in, U173_in, U174_in, U175_in, U176_in, U177_in, U178_in, U179_in, U180_in, U181_in, U182_in, U183_in, U184_in;
	wire signed [`WIDTH - 1:0] U176_in, U177_in, U178_in, U179_in, U180_in, U181_in, U182_in, U183_in, U184_in, U185_in, U186_in, U187_in, U188_in, U189_in, U190_in, U191_in;
	wire signed [`WIDTH - 1:0] U183_in, U184_in, U185_in, U186_in, U187_in, U188_in, U189_in, U190_in, U191_in, U192_in, U193_in, U194_in, U195_in, U196_in, U197_in, U198_in;
	wire signed [`WIDTH - 1:0] U190_in, U191_in, U192_in, U193_in, U194_in, U195_in, U196_in, U197_in, U198_in, U199_in, U200_in, U201_in, U202_in, U203_in, U204_in, U205_in;
	wire signed [`WIDTH - 1:0] U197_in, U198_in, U199_in, U200_in, U201_in, U202_in, U203_in, U204_in, U205_in, U206_in, U207_in, U208_in, U209_in, U210_in, U211_in, U212_in;
	wire signed [`WIDTH - 1:0] U204_in, U205_in, U206_in, U207_in, U208_in, U209_in, U210_in, U211_in, U212_in, U213_in, U214_in, U215_in, U216_in, U217_in, U218_in, U219_in;
	wire signed [`WIDTH - 1:0] U211_in, U212_in, U213_in, U214_in, U215_in, U216_in, U217_in, U218_in, U219_in, U220_in, U221_in, U222_in, U223_in, U224_in, U225_in, U226_in;
	wire signed [`WIDTH - 1:0] U218_in, U219_in, U220_in, U221_in, U222_in, U223_in, U224_in, U225_in, U226_in, U227_in, U228_in, U229_in, U230_in, U231_in, U232_in, U233_in;
	wire signed [`WIDTH - 1:0] U225_in, U226_in, U227_in, U228_in, U229_in, U230_in, U231_in, U232_in, U233_in, U234_in, U235_in, U236_in, U237_in, U238_in, U239_in, U240_in;
	wire signed [`WIDTH - 1:0] U232_in, U233_in, U234_in, U235_in, U236_in, U237_in, U238_in, U239_in, U240_in, U241_in, U242_in, U243_in, U244_in, U245_in, U246_in, U247_in;
	wire signed [`WIDTH - 1:0] U239_in, U240_in, U241_in, U242_in, U243_in, U244_in, U245_in, U246_in, U247_in, U248_in, U249_in, U250_in, U251_in, U252_in, U253_in, U254_in;
	wire signed [`WIDTH - 1:0] U246_in, U247_in, U248_in, U249_in, U250_in, U251_in, U252_in, U253_in, U254_in, U255_in, U256_in, U257_in, U258_in, U259_in, U260_in, U261_in;
	wire signed [`WIDTH - 1:0] U253_in, U254_in, U255_in, U256_in, U257_in, U258_in, U259_in, U260_in, U261_in, U262_in, U263_in, U264_in, U265_in, U266_in, U267_in, U268_in;
	wire signed [2 * `WIDTH - 1:0] Initial_X;
	output wire signed [2 * `WIDTH - 2:0] Y1_out, Y2_out, Y3_out, Y4_out, Y5_out, Y6_out, Y7_out, Y8_out, Y9_out, Y10_out, Y11_out, Y12_out, Y13_out, Y14_out, Y15_out, Y16_out;
	output wire signed [2 * `WIDTH - 2:0] Y8_out, Y9_out, Y10_out, Y11_out, Y12_out, Y13_out, Y14_out, Y15_out, Y16_out, Y17_out, Y18_out, Y19_out, Y20_out, Y21_out, Y22_out, Y23_out;
	output wire signed [2 * `WIDTH - 2:0] Y15_out, Y16_out, Y17_out, Y18_out, Y19_out, Y20_out, Y21_out, Y22_out, Y23_out, Y24_out, Y25_out, Y26_out, Y27_out, Y28_out, Y29_out, Y30_out;
	output wire signed [2 * `WIDTH - 2:0] Y22_out, Y23_out, Y24_out, Y25_out, Y26_out, Y27_out, Y28_out, Y29_out, Y30_out, Y31_out, Y32_out, Y33_out, Y34_out, Y35_out, Y36_out, Y37_out;
	output wire signed [2 * `WIDTH - 2:0] Y29_out, Y30_out, Y31_out, Y32_out, Y33_out, Y34_out, Y35_out, Y36_out, Y37_out, Y38_out, Y39_out, Y40_out, Y41_out, Y42_out, Y43_out, Y44_out;
	output wire signed [2 * `WIDTH - 2:0] Y36_out, Y37_out, Y38_out, Y39_out, Y40_out, Y41_out, Y42_out, Y43_out, Y44_out, Y45_out, Y46_out, Y47_out, Y48_out, Y49_out, Y50_out, Y51_out;
	output wire signed [2 * `WIDTH - 2:0] Y43_out, Y44_out, Y45_out, Y46_out, Y47_out, Y48_out, Y49_out, Y50_out, Y51_out, Y52_out, Y53_out, Y54_out, Y55_out, Y56_out, Y57_out, Y58_out;
	output wire signed [2 * `WIDTH - 2:0] Y50_out, Y51_out, Y52_out, Y53_out, Y54_out, Y55_out, Y56_out, Y57_out, Y58_out, Y59_out, Y60_out, Y61_out, Y62_out, Y63_out, Y64_out, Y65_out;
	output wire signed [2 * `WIDTH - 2:0] Y57_out, Y58_out, Y59_out, Y60_out, Y61_out, Y62_out, Y63_out, Y64_out, Y65_out, Y66_out, Y67_out, Y68_out, Y69_out, Y70_out, Y71_out, Y72_out;
	output wire signed [2 * `WIDTH - 2:0] Y64_out, Y65_out, Y66_out, Y67_out, Y68_out, Y69_out, Y70_out, Y71_out, Y72_out, Y73_out, Y74_out, Y75_out, Y76_out, Y77_out, Y78_out, Y79_out;
	output wire signed [2 * `WIDTH - 2:0] Y71_out, Y72_out, Y73_out, Y74_out, Y75_out, Y76_out, Y77_out, Y78_out, Y79_out, Y80_out, Y81_out, Y82_out, Y83_out, Y84_out, Y85_out, Y86_out;
	output wire signed [2 * `WIDTH - 2:0] Y78_out, Y79_out, Y80_out, Y81_out, Y82_out, Y83_out, Y84_out, Y85_out, Y86_out, Y87_out, Y88_out, Y89_out, Y90_out, Y91_out, Y92_out, Y93_out;
	output wire signed [2 * `WIDTH - 2:0] Y85_out, Y86_out, Y87_out, Y88_out, Y89_out, Y90_out, Y91_out, Y92_out, Y93_out, Y94_out, Y95_out, Y96_out, Y97_out, Y98_out, Y99_out, Y100_out;
	output wire signed [2 * `WIDTH - 2:0] Y92_out, Y93_out, Y94_out, Y95_out, Y96_out, Y97_out, Y98_out, Y99_out, Y100_out, Y101_out, Y102_out, Y103_out, Y104_out, Y105_out, Y106_out, Y107_out;
	output wire signed [2 * `WIDTH - 2:0] Y99_out, Y100_out, Y101_out, Y102_out, Y103_out, Y104_out, Y105_out, Y106_out, Y107_out, Y108_out, Y109_out, Y110_out, Y111_out, Y112_out, Y113_out, Y114_out;
	output wire signed [2 * `WIDTH - 2:0] Y106_out, Y107_out, Y108_out, Y109_out, Y110_out, Y111_out, Y112_out, Y113_out, Y114_out, Y115_out, Y116_out, Y117_out, Y118_out, Y119_out, Y120_out, Y121_out;
	output wire signed [2 * `WIDTH - 2:0] Y113_out, Y114_out, Y115_out, Y116_out, Y117_out, Y118_out, Y119_out, Y120_out, Y121_out, Y122_out, Y123_out, Y124_out, Y125_out, Y126_out, Y127_out, Y128_out;
	output wire signed [2 * `WIDTH - 2:0] Y120_out, Y121_out, Y122_out, Y123_out, Y124_out, Y125_out, Y126_out, Y127_out, Y128_out, Y129_out, Y130_out, Y131_out, Y132_out, Y133_out, Y134_out, Y135_out;
	output wire signed [2 * `WIDTH - 2:0] Y127_out, Y128_out, Y129_out, Y130_out, Y131_out, Y132_out, Y133_out, Y134_out, Y135_out, Y136_out, Y137_out, Y138_out, Y139_out, Y140_out, Y141_out, Y142_out;
	output wire signed [2 * `WIDTH - 2:0] Y134_out, Y135_out, Y136_out, Y137_out, Y138_out, Y139_out, Y140_out, Y141_out, Y142_out, Y143_out, Y144_out, Y145_out, Y146_out, Y147_out, Y148_out, Y149_out;
	output wire signed [2 * `WIDTH - 2:0] Y141_out, Y142_out, Y143_out, Y144_out, Y145_out, Y146_out, Y147_out, Y148_out, Y149_out, Y150_out, Y151_out, Y152_out, Y153_out, Y154_out, Y155_out, Y156_out;
	output wire signed [2 * `WIDTH - 2:0] Y148_out, Y149_out, Y150_out, Y151_out, Y152_out, Y153_out, Y154_out, Y155_out, Y156_out, Y157_out, Y158_out, Y159_out, Y160_out, Y161_out, Y162_out, Y163_out;
	output wire signed [2 * `WIDTH - 2:0] Y155_out, Y156_out, Y157_out, Y158_out, Y159_out, Y160_out, Y161_out, Y162_out, Y163_out, Y164_out, Y165_out, Y166_out, Y167_out, Y168_out, Y169_out, Y170_out;
	output wire signed [2 * `WIDTH - 2:0] Y162_out, Y163_out, Y164_out, Y165_out, Y166_out, Y167_out, Y168_out, Y169_out, Y170_out, Y171_out, Y172_out, Y173_out, Y174_out, Y175_out, Y176_out, Y177_out;
	output wire signed [2 * `WIDTH - 2:0] Y169_out, Y170_out, Y171_out, Y172_out, Y173_out, Y174_out, Y175_out, Y176_out, Y177_out, Y178_out, Y179_out, Y180_out, Y181_out, Y182_out, Y183_out, Y184_out;
	output wire signed [2 * `WIDTH - 2:0] Y176_out, Y177_out, Y178_out, Y179_out, Y180_out, Y181_out, Y182_out, Y183_out, Y184_out, Y185_out, Y186_out, Y187_out, Y188_out, Y189_out, Y190_out, Y191_out;
	output wire signed [2 * `WIDTH - 2:0] Y183_out, Y184_out, Y185_out, Y186_out, Y187_out, Y188_out, Y189_out, Y190_out, Y191_out, Y192_out, Y193_out, Y194_out, Y195_out, Y196_out, Y197_out, Y198_out;
	output wire signed [2 * `WIDTH - 2:0] Y190_out, Y191_out, Y192_out, Y193_out, Y194_out, Y195_out, Y196_out, Y197_out, Y198_out, Y199_out, Y200_out, Y201_out, Y202_out, Y203_out, Y204_out, Y205_out;
	output wire signed [2 * `WIDTH - 2:0] Y197_out, Y198_out, Y199_out, Y200_out, Y201_out, Y202_out, Y203_out, Y204_out, Y205_out, Y206_out, Y207_out, Y208_out, Y209_out, Y210_out, Y211_out, Y212_out;
	output wire signed [2 * `WIDTH - 2:0] Y204_out, Y205_out, Y206_out, Y207_out, Y208_out, Y209_out, Y210_out, Y211_out, Y212_out, Y213_out, Y214_out, Y215_out, Y216_out, Y217_out, Y218_out, Y219_out;
	output wire signed [2 * `WIDTH - 2:0] Y211_out, Y212_out, Y213_out, Y214_out, Y215_out, Y216_out, Y217_out, Y218_out, Y219_out, Y220_out, Y221_out, Y222_out, Y223_out, Y224_out, Y225_out, Y226_out;
	output wire signed [2 * `WIDTH - 2:0] Y218_out, Y219_out, Y220_out, Y221_out, Y222_out, Y223_out, Y224_out, Y225_out, Y226_out, Y227_out, Y228_out, Y229_out, Y230_out, Y231_out, Y232_out, Y233_out;
	output wire signed [2 * `WIDTH - 2:0] Y225_out, Y226_out, Y227_out, Y228_out, Y229_out, Y230_out, Y231_out, Y232_out, Y233_out, Y234_out, Y235_out, Y236_out, Y237_out, Y238_out, Y239_out, Y240_out;
	output wire signed [2 * `WIDTH - 2:0] Y232_out, Y233_out, Y234_out, Y235_out, Y236_out, Y237_out, Y238_out, Y239_out, Y240_out, Y241_out, Y242_out, Y243_out, Y244_out, Y245_out, Y246_out, Y247_out;
	output wire signed [2 * `WIDTH - 2:0] Y239_out, Y240_out, Y241_out, Y242_out, Y243_out, Y244_out, Y245_out, Y246_out, Y247_out, Y248_out, Y249_out, Y250_out, Y251_out, Y252_out, Y253_out, Y254_out;
	output wire signed [2 * `WIDTH - 2:0] Y246_out, Y247_out, Y248_out, Y249_out, Y250_out, Y251_out, Y252_out, Y253_out, Y254_out, Y255_out, Y256_out, Y257_out, Y258_out, Y259_out, Y260_out, Y261_out;
	output wire signed [2 * `WIDTH - 2:0] Y253_out, Y254_out, Y255_out, Y256_out, Y257_out, Y258_out, Y259_out, Y260_out, Y261_out, Y262_out, Y263_out, Y264_out, Y265_out, Y266_out, Y267_out, Y268_out;

//Value type is {signed, 2^3, 2^2, 2^1, 2^0, 2^-1...}
assign A1 = `WIDTH'b0;
assign A2 = `WIDTH'b0;
assign A3 = `WIDTH'b0;
assign A4 = `WIDTH'b0;
assign A5 = `WIDTH'b000010000;
assign A6 = `WIDTH'b0;
assign A7 = `WIDTH'b0;
assign A8 = `WIDTH'b0;
assign A9 = `WIDTH'b0;

assign B1 = `WIDTH'b111110000;
assign B2 = `WIDTH'b111110000;
assign B3 = `WIDTH'b111110000;
assign B4 = `WIDTH'b111110000;
assign B5 = `WIDTH'b001000000;
assign B6 = `WIDTH'b111110000;
assign B7 = `WIDTH'b111110000;
assign B8 = `WIDTH'b111110000;
assign B9 = `WIDTH'b111110000;
 
assign U1_out = `WIDTH'b0;assign U2_out = `WIDTH'b0;assign U3_out = `WIDTH'b0;assign U4_out = `WIDTH'b0;assign U5_out = `WIDTH'b0;assign U6_out = `WIDTH'b0;assign U7_out = `WIDTH'b0;assign U8_out = `WIDTH'b0;
assign U9_out = `WIDTH'b0;assign U10_out = `WIDTH'b0;assign U11_out = `WIDTH'b0;assign U12_out = `WIDTH'b0;assign U13_out = `WIDTH'b0;assign U14_out = `WIDTH'b0;assign U15_out = `WIDTH'b0;assign U16_out = `WIDTH'b0;
assign U17_out = `WIDTH'b0;assign U18_out = `WIDTH'b0;assign U19_out = `WIDTH'b0;assign U20_out = `WIDTH'b0;assign U21_out = `WIDTH'b0;assign U22_out = `WIDTH'b0;assign U23_out = `WIDTH'b0;assign U24_out = `WIDTH'b0;
assign U25_out = `WIDTH'b0;assign U26_out = `WIDTH'b0;assign U27_out = `WIDTH'b0;assign U28_out = `WIDTH'b0;assign U29_out = `WIDTH'b0;assign U30_out = `WIDTH'b0;assign U31_out = `WIDTH'b0;assign U32_out = `WIDTH'b0;
assign U33_out = `WIDTH'b0;assign U34_out = `WIDTH'b0;assign U35_out = `WIDTH'b0;assign U36_out = `WIDTH'b0;assign U37_out = `WIDTH'b0;assign U38_out = `WIDTH'b0;assign U39_out = `WIDTH'b0;assign U40_out = `WIDTH'b0;
assign U41_out = `WIDTH'b0;assign U42_out = `WIDTH'b0;assign U43_out = `WIDTH'b0;assign U44_out = `WIDTH'b0;assign U45_out = `WIDTH'b0;assign U46_out = `WIDTH'b0;assign U47_out = `WIDTH'b0;assign U48_out = `WIDTH'b0;
assign U49_out = `WIDTH'b0;assign U50_out = `WIDTH'b0;assign U51_out = `WIDTH'b0;assign U52_out = `WIDTH'b0;assign U53_out = `WIDTH'b0;assign U54_out = `WIDTH'b0;assign U55_out = `WIDTH'b0;assign U56_out = `WIDTH'b0;
assign U57_out = `WIDTH'b0;assign U58_out = `WIDTH'b0;assign U59_out = `WIDTH'b0;assign U60_out = `WIDTH'b0;assign U61_out = `WIDTH'b0;assign U62_out = `WIDTH'b0;assign U63_out = `WIDTH'b0;assign U64_out = `WIDTH'b0;
assign U65_out = `WIDTH'b0;assign U66_out = `WIDTH'b0;assign U67_out = `WIDTH'b0;assign U68_out = `WIDTH'b0;assign U69_out = `WIDTH'b0;assign U70_out = `WIDTH'b0;assign U71_out = `WIDTH'b0;assign U72_out = `WIDTH'b0;
assign U73_out = `WIDTH'b0;assign U74_out = `WIDTH'b0;assign U75_out = `WIDTH'b0;assign U76_out = `WIDTH'b0;assign U77_out = `WIDTH'b0;assign U78_out = `WIDTH'b0;assign U79_out = `WIDTH'b0;assign U80_out = `WIDTH'b0;
assign U81_out = `WIDTH'b0;assign U82_out = `WIDTH'b0;assign U83_out = `WIDTH'b0;assign U84_out = `WIDTH'b0;assign U85_out = `WIDTH'b0;assign U86_out = `WIDTH'b0;assign U87_out = `WIDTH'b0;assign U88_out = `WIDTH'b0;
assign U89_out = `WIDTH'b0;assign U90_out = `WIDTH'b0;assign U91_out = `WIDTH'b0;assign U92_out = `WIDTH'b0;assign U93_out = `WIDTH'b0;assign U94_out = `WIDTH'b0;assign U95_out = `WIDTH'b0;assign U96_out = `WIDTH'b0;
assign U97_out = `WIDTH'b0;assign U98_out = `WIDTH'b0;assign U99_out = `WIDTH'b0;assign U100_out = `WIDTH'b0;assign U101_out = `WIDTH'b0;assign U102_out = `WIDTH'b0;assign U103_out = `WIDTH'b0;assign U104_out = `WIDTH'b0;
assign U105_out = `WIDTH'b0;assign U106_out = `WIDTH'b0;assign U107_out = `WIDTH'b0;assign U108_out = `WIDTH'b0;assign U109_out = `WIDTH'b0;assign U110_out = `WIDTH'b0;assign U111_out = `WIDTH'b0;assign U112_out = `WIDTH'b0;
assign U113_out = `WIDTH'b0;assign U114_out = `WIDTH'b0;assign U115_out = `WIDTH'b0;assign U116_out = `WIDTH'b0;assign U117_out = `WIDTH'b0;assign U118_out = `WIDTH'b0;assign U119_out = `WIDTH'b0;assign U120_out = `WIDTH'b0;
assign U121_out = `WIDTH'b0;assign U122_out = `WIDTH'b0;assign U123_out = `WIDTH'b0;assign U124_out = `WIDTH'b0;assign U125_out = `WIDTH'b0;assign U126_out = `WIDTH'b0;assign U127_out = `WIDTH'b0;assign U128_out = `WIDTH'b0;
assign U129_out = `WIDTH'b0;assign U130_out = `WIDTH'b0;assign U131_out = `WIDTH'b0;assign U132_out = `WIDTH'b0;assign U133_out = `WIDTH'b0;assign U134_out = `WIDTH'b0;assign U135_out = `WIDTH'b0;assign U136_out = `WIDTH'b0;
assign U137_out = `WIDTH'b0;assign U138_out = `WIDTH'b0;assign U139_out = `WIDTH'b0;assign U140_out = `WIDTH'b0;assign U141_out = `WIDTH'b0;assign U142_out = `WIDTH'b0;assign U143_out = `WIDTH'b0;assign U144_out = `WIDTH'b0;
assign U145_out = `WIDTH'b0;assign U146_out = `WIDTH'b0;assign U147_out = `WIDTH'b0;assign U148_out = `WIDTH'b0;assign U149_out = `WIDTH'b0;assign U150_out = `WIDTH'b0;assign U151_out = `WIDTH'b0;assign U152_out = `WIDTH'b0;
assign U153_out = `WIDTH'b0;assign U154_out = `WIDTH'b0;assign U155_out = `WIDTH'b0;assign U156_out = `WIDTH'b0;assign U157_out = `WIDTH'b0;assign U158_out = `WIDTH'b0;assign U159_out = `WIDTH'b0;assign U160_out = `WIDTH'b0;
assign U161_out = `WIDTH'b0;assign U162_out = `WIDTH'b0;assign U163_out = `WIDTH'b0;assign U164_out = `WIDTH'b0;assign U165_out = `WIDTH'b0;assign U166_out = `WIDTH'b0;assign U167_out = `WIDTH'b0;assign U168_out = `WIDTH'b0;
assign U169_out = `WIDTH'b0;assign U170_out = `WIDTH'b0;assign U171_out = `WIDTH'b0;assign U172_out = `WIDTH'b0;assign U173_out = `WIDTH'b0;assign U174_out = `WIDTH'b0;assign U175_out = `WIDTH'b0;assign U176_out = `WIDTH'b0;
assign U177_out = `WIDTH'b0;assign U178_out = `WIDTH'b0;assign U179_out = `WIDTH'b0;assign U180_out = `WIDTH'b0;assign U181_out = `WIDTH'b0;assign U182_out = `WIDTH'b0;assign U183_out = `WIDTH'b0;assign U184_out = `WIDTH'b0;
assign U185_out = `WIDTH'b0;assign U186_out = `WIDTH'b0;assign U187_out = `WIDTH'b0;assign U188_out = `WIDTH'b0;assign U189_out = `WIDTH'b0;assign U190_out = `WIDTH'b0;assign U191_out = `WIDTH'b0;assign U192_out = `WIDTH'b0;
assign U193_out = `WIDTH'b0;assign U194_out = `WIDTH'b0;assign U195_out = `WIDTH'b0;assign U196_out = `WIDTH'b0;assign U197_out = `WIDTH'b0;assign U198_out = `WIDTH'b0;assign U199_out = `WIDTH'b0;assign U200_out = `WIDTH'b0;
assign U201_out = `WIDTH'b0;assign U202_out = `WIDTH'b0;assign U203_out = `WIDTH'b0;assign U204_out = `WIDTH'b0;assign U205_out = `WIDTH'b0;assign U206_out = `WIDTH'b0;assign U207_out = `WIDTH'b0;assign U208_out = `WIDTH'b0;
assign U209_out = `WIDTH'b0;assign U210_out = `WIDTH'b0;assign U211_out = `WIDTH'b0;assign U212_out = `WIDTH'b0;assign U213_out = `WIDTH'b0;assign U214_out = `WIDTH'b0;assign U215_out = `WIDTH'b0;assign U216_out = `WIDTH'b0;
assign U217_out = `WIDTH'b0;assign U218_out = `WIDTH'b0;assign U219_out = `WIDTH'b0;assign U220_out = `WIDTH'b0;assign U221_out = `WIDTH'b0;assign U222_out = `WIDTH'b0;assign U223_out = `WIDTH'b0;assign U224_out = `WIDTH'b0;
assign U225_out = `WIDTH'b0;assign U226_out = `WIDTH'b0;assign U227_out = `WIDTH'b0;assign U228_out = `WIDTH'b0;assign U229_out = `WIDTH'b0;assign U230_out = `WIDTH'b0;assign U231_out = `WIDTH'b0;assign U232_out = `WIDTH'b0;
assign U233_out = `WIDTH'b0;assign U234_out = `WIDTH'b0;assign U235_out = `WIDTH'b0;assign U236_out = `WIDTH'b0;assign U237_out = `WIDTH'b0;assign U238_out = `WIDTH'b0;assign U239_out = `WIDTH'b0;assign U240_out = `WIDTH'b0;
assign U241_out = `WIDTH'b0;assign U242_out = `WIDTH'b0;assign U243_out = `WIDTH'b0;assign U244_out = `WIDTH'b0;assign U245_out = `WIDTH'b0;assign U246_out = `WIDTH'b0;assign U247_out = `WIDTH'b0;assign U248_out = `WIDTH'b0;
assign U249_out = `WIDTH'b0;assign U250_out = `WIDTH'b0;assign U251_out = `WIDTH'b0;assign U252_out = `WIDTH'b0;assign U253_out = `WIDTH'b0;assign U254_out = `WIDTH'b0;assign U255_out = `WIDTH'b0;assign U256_out = `WIDTH'b0;


assign I = `WIDTH'b110110000;

assign Initial_X = {(2 * `WIDTH){1'b0}};

fourbyfour u1(

.clk(clk),

.A1(A1[`WIDTH - 1:0]),
.A2(A2[`WIDTH - 1:0]),
.A3(A3[`WIDTH - 1:0]),
.A4(A4[`WIDTH - 1:0]),
.A5(A5[`WIDTH - 1:0]),
.A6(A6[`WIDTH - 1:0]),
.A7(A7[`WIDTH - 1:0]),
.A8(A8[`WIDTH - 1:0]),
.A9(A9[`WIDTH - 1:0]),

.B1(B1[`WIDTH - 1:0]),
.B2(B2[`WIDTH - 1:0]),
.B3(B3[`WIDTH - 1:0]),
.B4(B4[`WIDTH - 1:0]),
.B5(B5[`WIDTH - 1:0]),
.B6(B6[`WIDTH - 1:0]),
.B7(B7[`WIDTH - 1:0]),
.B8(B8[`WIDTH - 1:0]),
.B9(B9[`WIDTH - 1:0]),

.U1_in(U1_in[`WIDTH - 1:0]),
.U2_in(U2_in[`WIDTH - 1:0]),
.U3_in(U3_in[`WIDTH - 1:0]),
.U4_in(U4_in[`WIDTH - 1:0]),
.U5_in(U5_in[`WIDTH - 1:0]),
.U6_in(U6_in[`WIDTH - 1:0]),
.U7_in(U7_in[`WIDTH - 1:0]),
.U8_in(U8_in[`WIDTH - 1:0]),
.U9_in(U9_in[`WIDTH - 1:0]),
.U10_in(U10_in[`WIDTH - 1:0]),
.U11_in(U11_in[`WIDTH - 1:0]),
.U12_in(U12_in[`WIDTH - 1:0]),
.U13_in(U13_in[`WIDTH - 1:0]),
.U14_in(U14_in[`WIDTH - 1:0]),
.U15_in(U15_in[`WIDTH - 1:0]),
.U16_in(U16_in[`WIDTH - 1:0]),

.Y1_out(Y1_out[2 * `WIDTH - 1:0]),
.Y2_out(Y2_out[2 * `WIDTH - 1:0]),
.Y3_out(Y3_out[2 * `WIDTH - 1:0]),
.Y4_out(Y4_out[2 * `WIDTH - 1:0]),
.Y5_out(Y5_out[2 * `WIDTH - 1:0]),
.Y6_out(Y6_out[2 * `WIDTH - 1:0]),
.Y7_out(Y7_out[2 * `WIDTH - 1:0]),
.Y8_out(Y8_out[2 * `WIDTH - 1:0]),
.Y9_out(Y9_out[2 * `WIDTH - 1:0]),
.Y10_out(Y10_out[2 * `WIDTH - 1:0]),
.Y11_out(Y11_out[2 * `WIDTH - 1:0]),
.Y12_out(Y12_out[2 * `WIDTH - 1:0]),
.Y13_out(Y13_out[2 * `WIDTH - 1:0]),
.Y14_out(Y14_out[2 * `WIDTH - 1:0]),
.Y15_out(Y15_out[2 * `WIDTH - 1:0]),
.Y16_out(Y16_out[2 * `WIDTH - 1:0]),

.I(I[`WIDTH - 1:0]),

.Initial_X_in(Initial_X[2 * `WIDTH - 1:0])
);

endmodule
