// The CNN module takes in the clock and give out the output matrix. 

`define WIDTH 9
module CNN (
clk,

Y1_out, Y2_out, Y3_out, Y4_out, Y5_out, Y6_out, Y7_out, Y8_out, Y9_out, Y10_out, Y11_out, Y12_out, Y13_out, Y14_out, Y15_out, Y16_out,
Y17_out, Y18_out, Y19_out, Y20_out, Y21_out, Y22_out, Y23_out, Y24_out, Y25_out, Y26_out, Y27_out, Y28_out, Y29_out, Y30_out, Y31_out, Y32_out,
Y33_out, Y34_out, Y35_out, Y36_out, Y37_out, Y38_out, Y39_out, Y40_out, Y41_out, Y42_out, Y43_out, Y44_out, Y45_out, Y46_out, Y47_out, Y48_out,
Y49_out, Y50_out, Y51_out, Y52_out, Y53_out, Y54_out, Y55_out, Y56_out, Y57_out, Y58_out, Y59_out, Y60_out, Y61_out, Y62_out, Y63_out, Y64_out,
Y65_out, Y66_out, Y67_out, Y68_out, Y69_out, Y70_out, Y71_out, Y72_out, Y73_out, Y74_out, Y75_out, Y76_out, Y77_out, Y78_out, Y79_out, Y80_out,
Y81_out, Y82_out, Y83_out, Y84_out, Y85_out, Y86_out, Y87_out, Y88_out, Y89_out, Y90_out, Y91_out, Y92_out, Y93_out, Y94_out, Y95_out, Y96_out,
Y97_out, Y98_out, Y99_out, Y100_out, Y101_out, Y102_out, Y103_out, Y104_out, Y105_out, Y106_out, Y107_out, Y108_out, Y109_out, Y110_out, Y111_out, Y112_out,
Y113_out, Y114_out, Y115_out, Y116_out, Y117_out, Y118_out, Y119_out, Y120_out, Y121_out, Y122_out, Y123_out, Y124_out, Y125_out, Y126_out, Y127_out, Y128_out,
Y129_out, Y130_out, Y131_out, Y132_out, Y133_out, Y134_out, Y135_out, Y136_out, Y137_out, Y138_out, Y139_out, Y140_out, Y141_out, Y142_out, Y143_out, Y144_out,
Y145_out, Y146_out, Y147_out, Y148_out, Y149_out, Y150_out, Y151_out, Y152_out, Y153_out, Y154_out, Y155_out, Y156_out, Y157_out, Y158_out, Y159_out, Y160_out,
Y161_out, Y162_out, Y163_out, Y164_out, Y165_out, Y166_out, Y167_out, Y168_out, Y169_out, Y170_out, Y171_out, Y172_out, Y173_out, Y174_out, Y175_out, Y176_out,
Y177_out, Y178_out, Y179_out, Y180_out, Y181_out, Y182_out, Y183_out, Y184_out, Y185_out, Y186_out, Y187_out, Y188_out, Y189_out, Y190_out, Y191_out, Y192_out,
Y193_out, Y194_out, Y195_out, Y196_out, Y197_out, Y198_out, Y199_out, Y200_out, Y201_out, Y202_out, Y203_out, Y204_out, Y205_out, Y206_out, Y207_out, Y208_out,
Y209_out, Y210_out, Y211_out, Y212_out, Y213_out, Y214_out, Y215_out, Y216_out, Y217_out, Y218_out, Y219_out, Y220_out, Y221_out, Y222_out, Y223_out, Y224_out,
Y225_out, Y226_out, Y227_out, Y228_out, Y229_out, Y230_out, Y231_out, Y232_out, Y233_out, Y234_out, Y235_out, Y236_out, Y237_out, Y238_out, Y239_out, Y240_out,
Y241_out, Y242_out, Y243_out, Y244_out, Y245_out, Y246_out, Y247_out, Y248_out, Y249_out, Y250_out, Y251_out, Y252_out, Y253_out, Y254_out, Y255_out, Y256_out

  );

// This module initializes all the inputs and gives it to the sixteenbysixteen module.
// It can similaly be given to onebyone or fourbyfour modules with respective lengths.
	input wire clk;
	wire signed [`WIDTH - 1:0] A1, A2, A3, A4, A5, A6, A7, A8, A9;
	wire signed [`WIDTH - 1:0] B1, B2, B3, B4, B5, B6, B7, B8, B9;
	wire signed [`WIDTH - 1:0] I;
	wire signed [`WIDTH - 1:0] U1_in, U2_in, U3_in, U4_in, U5_in, U6_in, U7_in, U8_in, U9_in, U10_in, U11_in, U12_in, U13_in, U14_in, U15_in, U16_in;
	wire signed [`WIDTH - 1:0] U17_in, U18_in, U19_in, U20_in, U21_in, U22_in, U23_in, U24_in, U25_in, U26_in, U27_in, U28_in, U29_in, U30_in, U31_in, U32_in;
	wire signed [`WIDTH - 1:0] U33_in, U34_in, U35_in, U36_in, U37_in, U38_in, U39_in, U40_in, U41_in, U42_in, U43_in, U44_in, U45_in, U46_in, U47_in, U48_in;
	wire signed [`WIDTH - 1:0] U49_in, U50_in, U51_in, U52_in, U53_in, U54_in, U55_in, U56_in, U57_in, U58_in, U59_in, U60_in, U61_in, U62_in, U63_in, U64_in;
	wire signed [`WIDTH - 1:0] U65_in, U66_in, U67_in, U68_in, U69_in, U70_in, U71_in, U72_in, U73_in, U74_in, U75_in, U76_in, U77_in, U78_in, U79_in, U80_in;
	wire signed [`WIDTH - 1:0] U81_in, U82_in, U83_in, U84_in, U85_in, U86_in, U87_in, U88_in, U89_in, U90_in, U91_in, U92_in, U93_in, U94_in, U95_in, U96_in;
	wire signed [`WIDTH - 1:0] U97_in, U98_in, U99_in, U100_in, U101_in, U102_in, U103_in, U104_in, U105_in, U106_in, U107_in, U108_in, U109_in, U110_in, U111_in, U112_in;
	wire signed [`WIDTH - 1:0] U113_in, U114_in, U115_in, U116_in, U117_in, U118_in, U119_in, U120_in, U121_in, U122_in, U123_in, U124_in, U125_in, U126_in, U127_in, U128_in;
	wire signed [`WIDTH - 1:0] U129_in, U130_in, U131_in, U132_in, U133_in, U134_in, U135_in, U136_in, U137_in, U138_in, U139_in, U140_in, U141_in, U142_in, U143_in, U144_in;
	wire signed [`WIDTH - 1:0] U145_in, U146_in, U147_in, U148_in, U149_in, U150_in, U151_in, U152_in, U153_in, U154_in, U155_in, U156_in, U157_in, U158_in, U159_in, U160_in;
	wire signed [`WIDTH - 1:0] U161_in, U162_in, U163_in, U164_in, U165_in, U166_in, U167_in, U168_in, U169_in, U170_in, U171_in, U172_in, U173_in, U174_in, U175_in, U176_in;
	wire signed [`WIDTH - 1:0] U177_in, U178_in, U179_in, U180_in, U181_in, U182_in, U183_in, U184_in, U185_in, U186_in, U187_in, U188_in, U189_in, U190_in, U191_in, U192_in;
	wire signed [`WIDTH - 1:0] U193_in, U194_in, U195_in, U196_in, U197_in, U198_in, U199_in, U200_in, U201_in, U202_in, U203_in, U204_in, U205_in, U206_in, U207_in, U208_in;
	wire signed [`WIDTH - 1:0] U209_in, U210_in, U211_in, U212_in, U213_in, U214_in, U215_in, U216_in, U217_in, U218_in, U219_in, U220_in, U221_in, U222_in, U223_in, U224_in;
	wire signed [`WIDTH - 1:0] U225_in, U226_in, U227_in, U228_in, U229_in, U230_in, U231_in, U232_in, U233_in, U234_in, U235_in, U236_in, U237_in, U238_in, U239_in, U240_in;
	wire signed [`WIDTH - 1:0] U241_in, U242_in, U243_in, U244_in, U245_in, U246_in, U247_in, U248_in, U249_in, U250_in, U251_in, U252_in, U253_in, U254_in, U255_in, U256_in;

	wire signed [2 * `WIDTH - 1:0] Initial_X;
	output wire signed [2 * `WIDTH - 1:0] Y1_out, Y2_out, Y3_out, Y4_out, Y5_out, Y6_out, Y7_out, Y8_out, Y9_out, Y10_out, Y11_out, Y12_out, Y13_out, Y14_out, Y15_out, Y16_out;
	output wire signed [2 * `WIDTH - 1:0] Y17_out, Y18_out, Y19_out, Y20_out, Y21_out, Y22_out, Y23_out, Y24_out, Y25_out, Y26_out, Y27_out, Y28_out, Y29_out, Y30_out, Y31_out, Y32_out;
	output wire signed [2 * `WIDTH - 1:0] Y33_out, Y34_out, Y35_out, Y36_out, Y37_out, Y38_out, Y39_out, Y40_out, Y41_out, Y42_out, Y43_out, Y44_out, Y45_out, Y46_out, Y47_out, Y48_out;
	output wire signed [2 * `WIDTH - 1:0] Y49_out, Y50_out, Y51_out, Y52_out, Y53_out, Y54_out, Y55_out, Y56_out, Y57_out, Y58_out, Y59_out, Y60_out, Y61_out, Y62_out, Y63_out, Y64_out;
	output wire signed [2 * `WIDTH - 1:0] Y65_out, Y66_out, Y67_out, Y68_out, Y69_out, Y70_out, Y71_out, Y72_out, Y73_out, Y74_out, Y75_out, Y76_out, Y77_out, Y78_out, Y79_out, Y80_out;
	output wire signed [2 * `WIDTH - 1:0] Y81_out, Y82_out, Y83_out, Y84_out, Y85_out, Y86_out, Y87_out, Y88_out, Y89_out, Y90_out, Y91_out, Y92_out, Y93_out, Y94_out, Y95_out, Y96_out;
	output wire signed [2 * `WIDTH - 1:0] Y97_out, Y98_out, Y99_out, Y100_out, Y101_out, Y102_out, Y103_out, Y104_out, Y105_out, Y106_out, Y107_out, Y108_out, Y109_out, Y110_out, Y111_out, Y112_out;
	output wire signed [2 * `WIDTH - 1:0] Y113_out, Y114_out, Y115_out, Y116_out, Y117_out, Y118_out, Y119_out, Y120_out, Y121_out, Y122_out, Y123_out, Y124_out, Y125_out, Y126_out, Y127_out, Y128_out;
	output wire signed [2 * `WIDTH - 1:0] Y129_out, Y130_out, Y131_out, Y132_out, Y133_out, Y134_out, Y135_out, Y136_out, Y137_out, Y138_out, Y139_out, Y140_out, Y141_out, Y142_out, Y143_out, Y144_out;
	output wire signed [2 * `WIDTH - 1:0] Y145_out, Y146_out, Y147_out, Y148_out, Y149_out, Y150_out, Y151_out, Y152_out, Y153_out, Y154_out, Y155_out, Y156_out, Y157_out, Y158_out, Y159_out, Y160_out;
	output wire signed [2 * `WIDTH - 1:0] Y161_out, Y162_out, Y163_out, Y164_out, Y165_out, Y166_out, Y167_out, Y168_out, Y169_out, Y170_out, Y171_out, Y172_out, Y173_out, Y174_out, Y175_out, Y176_out;
	output wire signed [2 * `WIDTH - 1:0] Y177_out, Y178_out, Y179_out, Y180_out, Y181_out, Y182_out, Y183_out, Y184_out, Y185_out, Y186_out, Y187_out, Y188_out, Y189_out, Y190_out, Y191_out, Y192_out;
	output wire signed [2 * `WIDTH - 1:0] Y193_out, Y194_out, Y195_out, Y196_out, Y197_out, Y198_out, Y199_out, Y200_out, Y201_out, Y202_out, Y203_out, Y204_out, Y205_out, Y206_out, Y207_out, Y208_out;
	output wire signed [2 * `WIDTH - 1:0] Y209_out, Y210_out, Y211_out, Y212_out, Y213_out, Y214_out, Y215_out, Y216_out, Y217_out, Y218_out, Y219_out, Y220_out, Y221_out, Y222_out, Y223_out, Y224_out;
	output wire signed [2 * `WIDTH - 1:0] Y225_out, Y226_out, Y227_out, Y228_out, Y229_out, Y230_out, Y231_out, Y232_out, Y233_out, Y234_out, Y235_out, Y236_out, Y237_out, Y238_out, Y239_out, Y240_out;
	output wire signed [2 * `WIDTH - 1:0] Y241_out, Y242_out, Y243_out, Y244_out, Y245_out, Y246_out, Y247_out, Y248_out, Y249_out, Y250_out, Y251_out, Y252_out, Y253_out, Y254_out, Y255_out, Y256_out;

//Value type is {signed, 2^3, 2^2, 2^1, 2^0, 2^-1...}
assign A1 = `WIDTH'b0;
assign A2 = `WIDTH'b0;
assign A3 = `WIDTH'b0;
assign A4 = `WIDTH'b0;
assign A5 = `WIDTH'b000010000;
assign A6 = `WIDTH'b0;
assign A7 = `WIDTH'b0;
assign A8 = `WIDTH'b0;
assign A9 = `WIDTH'b0;

assign B1 = `WIDTH'b111110000;
assign B2 = `WIDTH'b111110000;
assign B3 = `WIDTH'b111110000;
assign B4 = `WIDTH'b111110000;
assign B5 = `WIDTH'b001000000;
assign B6 = `WIDTH'b111110000;
assign B7 = `WIDTH'b111110000;
assign B8 = `WIDTH'b111110000;
assign B9 = `WIDTH'b111110000;
 
assign U1_in = `WIDTH'b0;assign U2_in = `WIDTH'b0;assign U3_in = `WIDTH'b0;assign U4_in = `WIDTH'b0;assign U5_in = `WIDTH'b0;assign U6_in = `WIDTH'b0;assign U7_in = `WIDTH'b0;assign U8_in = `WIDTH'b0;
assign U9_in = `WIDTH'b0;assign U10_in = `WIDTH'b0;assign U11_in = `WIDTH'b0;assign U12_in = `WIDTH'b0;assign U13_in = `WIDTH'b0;assign U14_in = `WIDTH'b0;assign U15_in = `WIDTH'b0;assign U16_in = `WIDTH'b0;
assign U17_in = `WIDTH'b0;assign U18_in = `WIDTH'b0;assign U19_in = `WIDTH'b0;assign U20_in = `WIDTH'b0;assign U21_in = `WIDTH'b0;assign U22_in = `WIDTH'b0;assign U23_in = `WIDTH'b0;assign U24_in = `WIDTH'b0;
assign U25_in = `WIDTH'b0;assign U26_in = `WIDTH'b0;assign U27_in = `WIDTH'b0;assign U28_in = `WIDTH'b0;assign U29_in = `WIDTH'b0;assign U30_in = `WIDTH'b0;assign U31_in = `WIDTH'b0;assign U32_in = `WIDTH'b0;
assign U33_in = `WIDTH'b0;assign U34_in = `WIDTH'b0;assign U35_in = `WIDTH'b0;assign U36_in = `WIDTH'b0;assign U37_in = `WIDTH'b0;assign U38_in = `WIDTH'b0;assign U39_in = `WIDTH'b0;assign U40_in = `WIDTH'b0;
assign U41_in = `WIDTH'b0;assign U42_in = `WIDTH'b0;assign U43_in = `WIDTH'b0;assign U44_in = `WIDTH'b0;assign U45_in = `WIDTH'b0;assign U46_in = `WIDTH'b0;assign U47_in = `WIDTH'b0;assign U48_in = `WIDTH'b0;
assign U49_in = `WIDTH'b0;assign U50_in = `WIDTH'b0;assign U51_in = `WIDTH'b0;assign U52_in = `WIDTH'b0;assign U53_in = `WIDTH'b0;assign U54_in = `WIDTH'b0;assign U55_in = `WIDTH'b0;assign U56_in = `WIDTH'b0;
assign U57_in = `WIDTH'b0;assign U58_in = `WIDTH'b0;assign U59_in = `WIDTH'b0;assign U60_in = `WIDTH'b0;assign U61_in = `WIDTH'b0;assign U62_in = `WIDTH'b0;assign U63_in = `WIDTH'b0;assign U64_in = `WIDTH'b0;
assign U65_in = `WIDTH'b0;assign U66_in = `WIDTH'b0;assign U67_in = `WIDTH'b0;assign U68_in = `WIDTH'b0;assign U69_in = `WIDTH'b0;assign U70_in = `WIDTH'b0;assign U71_in = `WIDTH'b000010000;assign U72_in = `WIDTH'b000010000;
assign U73_in = `WIDTH'b000010000;assign U74_in = `WIDTH'b000010000;assign U75_in = `WIDTH'b0;assign U76_in = `WIDTH'b0;assign U77_in = `WIDTH'b0;assign U78_in = `WIDTH'b0;assign U79_in = `WIDTH'b0;assign U80_in = `WIDTH'b0;
assign U81_in = `WIDTH'b0;assign U82_in = `WIDTH'b0;assign U83_in = `WIDTH'b0;assign U84_in = `WIDTH'b0;assign U85_in = `WIDTH'b0;assign U86_in = `WIDTH'b0;assign U87_in = `WIDTH'b000010000;assign U88_in = `WIDTH'b000010000;
assign U89_in = `WIDTH'b000010000;assign U90_in = `WIDTH'b000010000;assign U91_in = `WIDTH'b0;assign U92_in = `WIDTH'b0;assign U93_in = `WIDTH'b0;assign U94_in = `WIDTH'b0;assign U95_in = `WIDTH'b0;assign U96_in = `WIDTH'b0;
assign U97_in = `WIDTH'b0;assign U98_in = `WIDTH'b0;assign U99_in = `WIDTH'b0;assign U100_in = `WIDTH'b0;assign U101_in = `WIDTH'b0;assign U102_in = `WIDTH'b0;assign U103_in = `WIDTH'b000010000;assign U104_in = `WIDTH'b000010000;
assign U105_in = `WIDTH'b000010000;assign U106_in = `WIDTH'b000010000;assign U107_in = `WIDTH'b0;assign U108_in = `WIDTH'b0;assign U109_in = `WIDTH'b0;assign U110_in = `WIDTH'b0;assign U111_in = `WIDTH'b0;assign U112_in = `WIDTH'b0;
assign U113_in = `WIDTH'b0;assign U114_in = `WIDTH'b0;assign U115_in = `WIDTH'b0;assign U116_in = `WIDTH'b0;assign U117_in = `WIDTH'b0;assign U118_in = `WIDTH'b0;assign U119_in = `WIDTH'b000010000;assign U120_in = `WIDTH'b000010000;
assign U121_in = `WIDTH'b000010000;assign U122_in = `WIDTH'b000010000;assign U123_in = `WIDTH'b0;assign U124_in = `WIDTH'b0;assign U125_in = `WIDTH'b0;assign U126_in = `WIDTH'b0;assign U127_in = `WIDTH'b0;assign U128_in = `WIDTH'b0;
assign U129_in = `WIDTH'b0;assign U130_in = `WIDTH'b0;assign U131_in = `WIDTH'b0;assign U132_in = `WIDTH'b0;assign U133_in = `WIDTH'b0;assign U134_in = `WIDTH'b0;assign U135_in = `WIDTH'b000010000;assign U136_in = `WIDTH'b000010000;
assign U137_in = `WIDTH'b000010000;assign U138_in = `WIDTH'b000010000;assign U139_in = `WIDTH'b0;assign U140_in = `WIDTH'b0;assign U141_in = `WIDTH'b0;assign U142_in = `WIDTH'b0;assign U143_in = `WIDTH'b0;assign U144_in = `WIDTH'b0;
assign U145_in = `WIDTH'b0;assign U146_in = `WIDTH'b0;assign U147_in = `WIDTH'b0;assign U148_in = `WIDTH'b0;assign U149_in = `WIDTH'b0;assign U150_in = `WIDTH'b0;assign U151_in = `WIDTH'b0;assign U152_in = `WIDTH'b0;
assign U153_in = `WIDTH'b0;assign U154_in = `WIDTH'b0;assign U155_in = `WIDTH'b0;assign U156_in = `WIDTH'b0;assign U157_in = `WIDTH'b0;assign U158_in = `WIDTH'b0;assign U159_in = `WIDTH'b0;assign U160_in = `WIDTH'b0;
assign U161_in = `WIDTH'b0;assign U162_in = `WIDTH'b0;assign U163_in = `WIDTH'b0;assign U164_in = `WIDTH'b0;assign U165_in = `WIDTH'b0;assign U166_in = `WIDTH'b0;assign U167_in = `WIDTH'b0;assign U168_in = `WIDTH'b0;
assign U169_in = `WIDTH'b0;assign U170_in = `WIDTH'b0;assign U171_in = `WIDTH'b0;assign U172_in = `WIDTH'b0;assign U173_in = `WIDTH'b0;assign U174_in = `WIDTH'b0;assign U175_in = `WIDTH'b0;assign U176_in = `WIDTH'b0;
assign U177_in = `WIDTH'b0;assign U178_in = `WIDTH'b0;assign U179_in = `WIDTH'b0;assign U180_in = `WIDTH'b0;assign U181_in = `WIDTH'b0;assign U182_in = `WIDTH'b0;assign U183_in = `WIDTH'b0;assign U184_in = `WIDTH'b0;
assign U185_in = `WIDTH'b0;assign U186_in = `WIDTH'b0;assign U187_in = `WIDTH'b0;assign U188_in = `WIDTH'b0;assign U189_in = `WIDTH'b0;assign U190_in = `WIDTH'b0;assign U191_in = `WIDTH'b0;assign U192_in = `WIDTH'b0;
assign U193_in = `WIDTH'b0;assign U194_in = `WIDTH'b0;assign U195_in = `WIDTH'b0;assign U196_in = `WIDTH'b0;assign U197_in = `WIDTH'b0;assign U198_in = `WIDTH'b0;assign U199_in = `WIDTH'b0;assign U200_in = `WIDTH'b0;
assign U201_in = `WIDTH'b0;assign U202_in = `WIDTH'b0;assign U203_in = `WIDTH'b0;assign U204_in = `WIDTH'b0;assign U205_in = `WIDTH'b0;assign U206_in = `WIDTH'b0;assign U207_in = `WIDTH'b0;assign U208_in = `WIDTH'b0;
assign U209_in = `WIDTH'b0;assign U210_in = `WIDTH'b0;assign U211_in = `WIDTH'b0;assign U212_in = `WIDTH'b0;assign U213_in = `WIDTH'b0;assign U214_in = `WIDTH'b0;assign U215_in = `WIDTH'b0;assign U216_in = `WIDTH'b0;
assign U217_in = `WIDTH'b0;assign U218_in = `WIDTH'b0;assign U219_in = `WIDTH'b0;assign U220_in = `WIDTH'b0;assign U221_in = `WIDTH'b0;assign U222_in = `WIDTH'b0;assign U223_in = `WIDTH'b0;assign U224_in = `WIDTH'b0;
assign U225_in = `WIDTH'b0;assign U226_in = `WIDTH'b0;assign U227_in = `WIDTH'b0;assign U228_in = `WIDTH'b0;assign U229_in = `WIDTH'b0;assign U230_in = `WIDTH'b0;assign U231_in = `WIDTH'b0;assign U232_in = `WIDTH'b0;
assign U233_in = `WIDTH'b0;assign U234_in = `WIDTH'b0;assign U235_in = `WIDTH'b0;assign U236_in = `WIDTH'b0;assign U237_in = `WIDTH'b0;assign U238_in = `WIDTH'b0;assign U239_in = `WIDTH'b0;assign U240_in = `WIDTH'b0;
assign U241_in = `WIDTH'b0;assign U242_in = `WIDTH'b0;assign U243_in = `WIDTH'b0;assign U244_in = `WIDTH'b0;assign U245_in = `WIDTH'b0;assign U246_in = `WIDTH'b0;assign U247_in = `WIDTH'b0;assign U248_in = `WIDTH'b0;
assign U249_in = `WIDTH'b0;assign U250_in = `WIDTH'b0;assign U251_in = `WIDTH'b0;assign U252_in = `WIDTH'b0;assign U253_in = `WIDTH'b0;assign U254_in = `WIDTH'b0;assign U255_in = `WIDTH'b0;assign U256_in = `WIDTH'b0;

assign I = `WIDTH'b110110000;

assign Initial_X = {(2 * `WIDTH){1'b0}};

sixteenbysixteen u1(

.clk(clk),

.A1(A1[`WIDTH - 1:0]),
.A2(A2[`WIDTH - 1:0]),
.A3(A3[`WIDTH - 1:0]),
.A4(A4[`WIDTH - 1:0]),
.A5(A5[`WIDTH - 1:0]),
.A6(A6[`WIDTH - 1:0]),
.A7(A7[`WIDTH - 1:0]),
.A8(A8[`WIDTH - 1:0]),
.A9(A9[`WIDTH - 1:0]),

.B1(B1[`WIDTH - 1:0]),
.B2(B2[`WIDTH - 1:0]),
.B3(B3[`WIDTH - 1:0]),
.B4(B4[`WIDTH - 1:0]),
.B5(B5[`WIDTH - 1:0]),
.B6(B6[`WIDTH - 1:0]),
.B7(B7[`WIDTH - 1:0]),
.B8(B8[`WIDTH - 1:0]),
.B9(B9[`WIDTH - 1:0]),

.U1_in(U1_in[`WIDTH - 1:0]),.U2_in(U2_in[`WIDTH - 1:0]),.U3_in(U3_in[`WIDTH - 1:0]),.U4_in(U4_in[`WIDTH - 1:0]),.U5_in(U5_in[`WIDTH - 1:0]),.U6_in(U6_in[`WIDTH - 1:0]),.U7_in(U7_in[`WIDTH - 1:0]),.U8_in(U8_in[`WIDTH - 1:0]),
.U9_in(U9_in[`WIDTH - 1:0]),.U10_in(U10_in[`WIDTH - 1:0]),.U11_in(U11_in[`WIDTH - 1:0]),.U12_in(U12_in[`WIDTH - 1:0]),.U13_in(U13_in[`WIDTH - 1:0]),.U14_in(U14_in[`WIDTH - 1:0]),.U15_in(U15_in[`WIDTH - 1:0]),.U16_in(U16_in[`WIDTH - 1:0]),
.U17_in(U17_in[`WIDTH - 1:0]),.U18_in(U18_in[`WIDTH - 1:0]),.U19_in(U19_in[`WIDTH - 1:0]),.U20_in(U20_in[`WIDTH - 1:0]),.U21_in(U21_in[`WIDTH - 1:0]),.U22_in(U22_in[`WIDTH - 1:0]),.U23_in(U23_in[`WIDTH - 1:0]),.U24_in(U24_in[`WIDTH - 1:0]),
.U25_in(U25_in[`WIDTH - 1:0]),.U26_in(U26_in[`WIDTH - 1:0]),.U27_in(U27_in[`WIDTH - 1:0]),.U28_in(U28_in[`WIDTH - 1:0]),.U29_in(U29_in[`WIDTH - 1:0]),.U30_in(U30_in[`WIDTH - 1:0]),.U31_in(U31_in[`WIDTH - 1:0]),.U32_in(U32_in[`WIDTH - 1:0]),
.U33_in(U33_in[`WIDTH - 1:0]),.U34_in(U34_in[`WIDTH - 1:0]),.U35_in(U35_in[`WIDTH - 1:0]),.U36_in(U36_in[`WIDTH - 1:0]),.U37_in(U37_in[`WIDTH - 1:0]),.U38_in(U38_in[`WIDTH - 1:0]),.U39_in(U39_in[`WIDTH - 1:0]),.U40_in(U40_in[`WIDTH - 1:0]),
.U41_in(U41_in[`WIDTH - 1:0]),.U42_in(U42_in[`WIDTH - 1:0]),.U43_in(U43_in[`WIDTH - 1:0]),.U44_in(U44_in[`WIDTH - 1:0]),.U45_in(U45_in[`WIDTH - 1:0]),.U46_in(U46_in[`WIDTH - 1:0]),.U47_in(U47_in[`WIDTH - 1:0]),.U48_in(U48_in[`WIDTH - 1:0]),
.U49_in(U49_in[`WIDTH - 1:0]),.U50_in(U50_in[`WIDTH - 1:0]),.U51_in(U51_in[`WIDTH - 1:0]),.U52_in(U52_in[`WIDTH - 1:0]),.U53_in(U53_in[`WIDTH - 1:0]),.U54_in(U54_in[`WIDTH - 1:0]),.U55_in(U55_in[`WIDTH - 1:0]),.U56_in(U56_in[`WIDTH - 1:0]),
.U57_in(U57_in[`WIDTH - 1:0]),.U58_in(U58_in[`WIDTH - 1:0]),.U59_in(U59_in[`WIDTH - 1:0]),.U60_in(U60_in[`WIDTH - 1:0]),.U61_in(U61_in[`WIDTH - 1:0]),.U62_in(U62_in[`WIDTH - 1:0]),.U63_in(U63_in[`WIDTH - 1:0]),.U64_in(U64_in[`WIDTH - 1:0]),
.U65_in(U65_in[`WIDTH - 1:0]),.U66_in(U66_in[`WIDTH - 1:0]),.U67_in(U67_in[`WIDTH - 1:0]),.U68_in(U68_in[`WIDTH - 1:0]),.U69_in(U69_in[`WIDTH - 1:0]),.U70_in(U70_in[`WIDTH - 1:0]),.U71_in(U71_in[`WIDTH - 1:0]),.U72_in(U72_in[`WIDTH - 1:0]),
.U73_in(U73_in[`WIDTH - 1:0]),.U74_in(U74_in[`WIDTH - 1:0]),.U75_in(U75_in[`WIDTH - 1:0]),.U76_in(U76_in[`WIDTH - 1:0]),.U77_in(U77_in[`WIDTH - 1:0]),.U78_in(U78_in[`WIDTH - 1:0]),.U79_in(U79_in[`WIDTH - 1:0]),.U80_in(U80_in[`WIDTH - 1:0]),
.U81_in(U81_in[`WIDTH - 1:0]),.U82_in(U82_in[`WIDTH - 1:0]),.U83_in(U83_in[`WIDTH - 1:0]),.U84_in(U84_in[`WIDTH - 1:0]),.U85_in(U85_in[`WIDTH - 1:0]),.U86_in(U86_in[`WIDTH - 1:0]),.U87_in(U87_in[`WIDTH - 1:0]),.U88_in(U88_in[`WIDTH - 1:0]),
.U89_in(U89_in[`WIDTH - 1:0]),.U90_in(U90_in[`WIDTH - 1:0]),.U91_in(U91_in[`WIDTH - 1:0]),.U92_in(U92_in[`WIDTH - 1:0]),.U93_in(U93_in[`WIDTH - 1:0]),.U94_in(U94_in[`WIDTH - 1:0]),.U95_in(U95_in[`WIDTH - 1:0]),.U96_in(U96_in[`WIDTH - 1:0]),
.U97_in(U97_in[`WIDTH - 1:0]),.U98_in(U98_in[`WIDTH - 1:0]),.U99_in(U99_in[`WIDTH - 1:0]),.U100_in(U100_in[`WIDTH - 1:0]),.U101_in(U101_in[`WIDTH - 1:0]),.U102_in(U102_in[`WIDTH - 1:0]),.U103_in(U103_in[`WIDTH - 1:0]),.U104_in(U104_in[`WIDTH - 1:0]),
.U105_in(U105_in[`WIDTH - 1:0]),.U106_in(U106_in[`WIDTH - 1:0]),.U107_in(U107_in[`WIDTH - 1:0]),.U108_in(U108_in[`WIDTH - 1:0]),.U109_in(U109_in[`WIDTH - 1:0]),.U110_in(U110_in[`WIDTH - 1:0]),.U111_in(U111_in[`WIDTH - 1:0]),.U112_in(U112_in[`WIDTH - 1:0]),
.U113_in(U113_in[`WIDTH - 1:0]),.U114_in(U114_in[`WIDTH - 1:0]),.U115_in(U115_in[`WIDTH - 1:0]),.U116_in(U116_in[`WIDTH - 1:0]),.U117_in(U117_in[`WIDTH - 1:0]),.U118_in(U118_in[`WIDTH - 1:0]),.U119_in(U119_in[`WIDTH - 1:0]),.U120_in(U120_in[`WIDTH - 1:0]),
.U121_in(U121_in[`WIDTH - 1:0]),.U122_in(U122_in[`WIDTH - 1:0]),.U123_in(U123_in[`WIDTH - 1:0]),.U124_in(U124_in[`WIDTH - 1:0]),.U125_in(U125_in[`WIDTH - 1:0]),.U126_in(U126_in[`WIDTH - 1:0]),.U127_in(U127_in[`WIDTH - 1:0]),.U128_in(U128_in[`WIDTH - 1:0]),
.U129_in(U129_in[`WIDTH - 1:0]),.U130_in(U130_in[`WIDTH - 1:0]),.U131_in(U131_in[`WIDTH - 1:0]),.U132_in(U132_in[`WIDTH - 1:0]),.U133_in(U133_in[`WIDTH - 1:0]),.U134_in(U134_in[`WIDTH - 1:0]),.U135_in(U135_in[`WIDTH - 1:0]),.U136_in(U136_in[`WIDTH - 1:0]),
.U137_in(U137_in[`WIDTH - 1:0]),.U138_in(U138_in[`WIDTH - 1:0]),.U139_in(U139_in[`WIDTH - 1:0]),.U140_in(U140_in[`WIDTH - 1:0]),.U141_in(U141_in[`WIDTH - 1:0]),.U142_in(U142_in[`WIDTH - 1:0]),.U143_in(U143_in[`WIDTH - 1:0]),.U144_in(U144_in[`WIDTH - 1:0]),
.U145_in(U145_in[`WIDTH - 1:0]),.U146_in(U146_in[`WIDTH - 1:0]),.U147_in(U147_in[`WIDTH - 1:0]),.U148_in(U148_in[`WIDTH - 1:0]),.U149_in(U149_in[`WIDTH - 1:0]),.U150_in(U150_in[`WIDTH - 1:0]),.U151_in(U151_in[`WIDTH - 1:0]),.U152_in(U152_in[`WIDTH - 1:0]),
.U153_in(U153_in[`WIDTH - 1:0]),.U154_in(U154_in[`WIDTH - 1:0]),.U155_in(U155_in[`WIDTH - 1:0]),.U156_in(U156_in[`WIDTH - 1:0]),.U157_in(U157_in[`WIDTH - 1:0]),.U158_in(U158_in[`WIDTH - 1:0]),.U159_in(U159_in[`WIDTH - 1:0]),.U160_in(U160_in[`WIDTH - 1:0]),
.U161_in(U161_in[`WIDTH - 1:0]),.U162_in(U162_in[`WIDTH - 1:0]),.U163_in(U163_in[`WIDTH - 1:0]),.U164_in(U164_in[`WIDTH - 1:0]),.U165_in(U165_in[`WIDTH - 1:0]),.U166_in(U166_in[`WIDTH - 1:0]),.U167_in(U167_in[`WIDTH - 1:0]),.U168_in(U168_in[`WIDTH - 1:0]),
.U169_in(U169_in[`WIDTH - 1:0]),.U170_in(U170_in[`WIDTH - 1:0]),.U171_in(U171_in[`WIDTH - 1:0]),.U172_in(U172_in[`WIDTH - 1:0]),.U173_in(U173_in[`WIDTH - 1:0]),.U174_in(U174_in[`WIDTH - 1:0]),.U175_in(U175_in[`WIDTH - 1:0]),.U176_in(U176_in[`WIDTH - 1:0]),
.U177_in(U177_in[`WIDTH - 1:0]),.U178_in(U178_in[`WIDTH - 1:0]),.U179_in(U179_in[`WIDTH - 1:0]),.U180_in(U180_in[`WIDTH - 1:0]),.U181_in(U181_in[`WIDTH - 1:0]),.U182_in(U182_in[`WIDTH - 1:0]),.U183_in(U183_in[`WIDTH - 1:0]),.U184_in(U184_in[`WIDTH - 1:0]),
.U185_in(U185_in[`WIDTH - 1:0]),.U186_in(U186_in[`WIDTH - 1:0]),.U187_in(U187_in[`WIDTH - 1:0]),.U188_in(U188_in[`WIDTH - 1:0]),.U189_in(U189_in[`WIDTH - 1:0]),.U190_in(U190_in[`WIDTH - 1:0]),.U191_in(U191_in[`WIDTH - 1:0]),.U192_in(U192_in[`WIDTH - 1:0]),
.U193_in(U193_in[`WIDTH - 1:0]),.U194_in(U194_in[`WIDTH - 1:0]),.U195_in(U195_in[`WIDTH - 1:0]),.U196_in(U196_in[`WIDTH - 1:0]),.U197_in(U197_in[`WIDTH - 1:0]),.U198_in(U198_in[`WIDTH - 1:0]),.U199_in(U199_in[`WIDTH - 1:0]),.U200_in(U200_in[`WIDTH - 1:0]),
.U201_in(U201_in[`WIDTH - 1:0]),.U202_in(U202_in[`WIDTH - 1:0]),.U203_in(U203_in[`WIDTH - 1:0]),.U204_in(U204_in[`WIDTH - 1:0]),.U205_in(U205_in[`WIDTH - 1:0]),.U206_in(U206_in[`WIDTH - 1:0]),.U207_in(U207_in[`WIDTH - 1:0]),.U208_in(U208_in[`WIDTH - 1:0]),
.U209_in(U209_in[`WIDTH - 1:0]),.U210_in(U210_in[`WIDTH - 1:0]),.U211_in(U211_in[`WIDTH - 1:0]),.U212_in(U212_in[`WIDTH - 1:0]),.U213_in(U213_in[`WIDTH - 1:0]),.U214_in(U214_in[`WIDTH - 1:0]),.U215_in(U215_in[`WIDTH - 1:0]),.U216_in(U216_in[`WIDTH - 1:0]),
.U217_in(U217_in[`WIDTH - 1:0]),.U218_in(U218_in[`WIDTH - 1:0]),.U219_in(U219_in[`WIDTH - 1:0]),.U220_in(U220_in[`WIDTH - 1:0]),.U221_in(U221_in[`WIDTH - 1:0]),.U222_in(U222_in[`WIDTH - 1:0]),.U223_in(U223_in[`WIDTH - 1:0]),.U224_in(U224_in[`WIDTH - 1:0]),
.U225_in(U225_in[`WIDTH - 1:0]),.U226_in(U226_in[`WIDTH - 1:0]),.U227_in(U227_in[`WIDTH - 1:0]),.U228_in(U228_in[`WIDTH - 1:0]),.U229_in(U229_in[`WIDTH - 1:0]),.U230_in(U230_in[`WIDTH - 1:0]),.U231_in(U231_in[`WIDTH - 1:0]),.U232_in(U232_in[`WIDTH - 1:0]),
.U233_in(U233_in[`WIDTH - 1:0]),.U234_in(U234_in[`WIDTH - 1:0]),.U235_in(U235_in[`WIDTH - 1:0]),.U236_in(U236_in[`WIDTH - 1:0]),.U237_in(U237_in[`WIDTH - 1:0]),.U238_in(U238_in[`WIDTH - 1:0]),.U239_in(U239_in[`WIDTH - 1:0]),.U240_in(U240_in[`WIDTH - 1:0]),
.U241_in(U241_in[`WIDTH - 1:0]),.U242_in(U242_in[`WIDTH - 1:0]),.U243_in(U243_in[`WIDTH - 1:0]),.U244_in(U244_in[`WIDTH - 1:0]),.U245_in(U245_in[`WIDTH - 1:0]),.U246_in(U246_in[`WIDTH - 1:0]),.U247_in(U247_in[`WIDTH - 1:0]),.U248_in(U248_in[`WIDTH - 1:0]),
.U249_in(U249_in[`WIDTH - 1:0]),.U250_in(U250_in[`WIDTH - 1:0]),.U251_in(U251_in[`WIDTH - 1:0]),.U252_in(U252_in[`WIDTH - 1:0]),.U253_in(U253_in[`WIDTH - 1:0]),.U254_in(U254_in[`WIDTH - 1:0]),.U255_in(U255_in[`WIDTH - 1:0]),.U256_in(U256_in[`WIDTH - 1:0]),

.Y1_out(Y1_out[2 * `WIDTH - 1:0]),.Y2_out(Y2_out[2 * `WIDTH - 1:0]),.Y3_out(Y3_out[2 * `WIDTH - 1:0]),.Y4_out(Y4_out[2 * `WIDTH - 1:0]),.Y5_out(Y5_out[2 * `WIDTH - 1:0]),.Y6_out(Y6_out[2 * `WIDTH - 1:0]),.Y7_out(Y7_out[2 * `WIDTH - 1:0]),.Y8_out(Y8_out[2 * `WIDTH - 1:0]),
.Y9_out(Y9_out[2 * `WIDTH - 1:0]),.Y10_out(Y10_out[2 * `WIDTH - 1:0]),.Y11_out(Y11_out[2 * `WIDTH - 1:0]),.Y12_out(Y12_out[2 * `WIDTH - 1:0]),.Y13_out(Y13_out[2 * `WIDTH - 1:0]),.Y14_out(Y14_out[2 * `WIDTH - 1:0]),.Y15_out(Y15_out[2 * `WIDTH - 1:0]),.Y16_out(Y16_out[2 * `WIDTH - 1:0]),
.Y17_out(Y17_out[2 * `WIDTH - 1:0]),.Y18_out(Y18_out[2 * `WIDTH - 1:0]),.Y19_out(Y19_out[2 * `WIDTH - 1:0]),.Y20_out(Y20_out[2 * `WIDTH - 1:0]),.Y21_out(Y21_out[2 * `WIDTH - 1:0]),.Y22_out(Y22_out[2 * `WIDTH - 1:0]),.Y23_out(Y23_out[2 * `WIDTH - 1:0]),.Y24_out(Y24_out[2 * `WIDTH - 1:0]),
.Y25_out(Y25_out[2 * `WIDTH - 1:0]),.Y26_out(Y26_out[2 * `WIDTH - 1:0]),.Y27_out(Y27_out[2 * `WIDTH - 1:0]),.Y28_out(Y28_out[2 * `WIDTH - 1:0]),.Y29_out(Y29_out[2 * `WIDTH - 1:0]),.Y30_out(Y30_out[2 * `WIDTH - 1:0]),.Y31_out(Y31_out[2 * `WIDTH - 1:0]),.Y32_out(Y32_out[2 * `WIDTH - 1:0]),
.Y33_out(Y33_out[2 * `WIDTH - 1:0]),.Y34_out(Y34_out[2 * `WIDTH - 1:0]),.Y35_out(Y35_out[2 * `WIDTH - 1:0]),.Y36_out(Y36_out[2 * `WIDTH - 1:0]),.Y37_out(Y37_out[2 * `WIDTH - 1:0]),.Y38_out(Y38_out[2 * `WIDTH - 1:0]),.Y39_out(Y39_out[2 * `WIDTH - 1:0]),.Y40_out(Y40_out[2 * `WIDTH - 1:0]),
.Y41_out(Y41_out[2 * `WIDTH - 1:0]),.Y42_out(Y42_out[2 * `WIDTH - 1:0]),.Y43_out(Y43_out[2 * `WIDTH - 1:0]),.Y44_out(Y44_out[2 * `WIDTH - 1:0]),.Y45_out(Y45_out[2 * `WIDTH - 1:0]),.Y46_out(Y46_out[2 * `WIDTH - 1:0]),.Y47_out(Y47_out[2 * `WIDTH - 1:0]),.Y48_out(Y48_out[2 * `WIDTH - 1:0]),
.Y49_out(Y49_out[2 * `WIDTH - 1:0]),.Y50_out(Y50_out[2 * `WIDTH - 1:0]),.Y51_out(Y51_out[2 * `WIDTH - 1:0]),.Y52_out(Y52_out[2 * `WIDTH - 1:0]),.Y53_out(Y53_out[2 * `WIDTH - 1:0]),.Y54_out(Y54_out[2 * `WIDTH - 1:0]),.Y55_out(Y55_out[2 * `WIDTH - 1:0]),.Y56_out(Y56_out[2 * `WIDTH - 1:0]),
.Y57_out(Y57_out[2 * `WIDTH - 1:0]),.Y58_out(Y58_out[2 * `WIDTH - 1:0]),.Y59_out(Y59_out[2 * `WIDTH - 1:0]),.Y60_out(Y60_out[2 * `WIDTH - 1:0]),.Y61_out(Y61_out[2 * `WIDTH - 1:0]),.Y62_out(Y62_out[2 * `WIDTH - 1:0]),.Y63_out(Y63_out[2 * `WIDTH - 1:0]),.Y64_out(Y64_out[2 * `WIDTH - 1:0]),
.Y65_out(Y65_out[2 * `WIDTH - 1:0]),.Y66_out(Y66_out[2 * `WIDTH - 1:0]),.Y67_out(Y67_out[2 * `WIDTH - 1:0]),.Y68_out(Y68_out[2 * `WIDTH - 1:0]),.Y69_out(Y69_out[2 * `WIDTH - 1:0]),.Y70_out(Y70_out[2 * `WIDTH - 1:0]),.Y71_out(Y71_out[2 * `WIDTH - 1:0]),.Y72_out(Y72_out[2 * `WIDTH - 1:0]),
.Y73_out(Y73_out[2 * `WIDTH - 1:0]),.Y74_out(Y74_out[2 * `WIDTH - 1:0]),.Y75_out(Y75_out[2 * `WIDTH - 1:0]),.Y76_out(Y76_out[2 * `WIDTH - 1:0]),.Y77_out(Y77_out[2 * `WIDTH - 1:0]),.Y78_out(Y78_out[2 * `WIDTH - 1:0]),.Y79_out(Y79_out[2 * `WIDTH - 1:0]),.Y80_out(Y80_out[2 * `WIDTH - 1:0]),
.Y81_out(Y81_out[2 * `WIDTH - 1:0]),.Y82_out(Y82_out[2 * `WIDTH - 1:0]),.Y83_out(Y83_out[2 * `WIDTH - 1:0]),.Y84_out(Y84_out[2 * `WIDTH - 1:0]),.Y85_out(Y85_out[2 * `WIDTH - 1:0]),.Y86_out(Y86_out[2 * `WIDTH - 1:0]),.Y87_out(Y87_out[2 * `WIDTH - 1:0]),.Y88_out(Y88_out[2 * `WIDTH - 1:0]),
.Y89_out(Y89_out[2 * `WIDTH - 1:0]),.Y90_out(Y90_out[2 * `WIDTH - 1:0]),.Y91_out(Y91_out[2 * `WIDTH - 1:0]),.Y92_out(Y92_out[2 * `WIDTH - 1:0]),.Y93_out(Y93_out[2 * `WIDTH - 1:0]),.Y94_out(Y94_out[2 * `WIDTH - 1:0]),.Y95_out(Y95_out[2 * `WIDTH - 1:0]),.Y96_out(Y96_out[2 * `WIDTH - 1:0]),
.Y97_out(Y97_out[2 * `WIDTH - 1:0]),.Y98_out(Y98_out[2 * `WIDTH - 1:0]),.Y99_out(Y99_out[2 * `WIDTH - 1:0]),.Y100_out(Y100_out[2 * `WIDTH - 1:0]),.Y101_out(Y101_out[2 * `WIDTH - 1:0]),.Y102_out(Y102_out[2 * `WIDTH - 1:0]),.Y103_out(Y103_out[2 * `WIDTH - 1:0]),.Y104_out(Y104_out[2 * `WIDTH - 1:0]),
.Y105_out(Y105_out[2 * `WIDTH - 1:0]),.Y106_out(Y106_out[2 * `WIDTH - 1:0]),.Y107_out(Y107_out[2 * `WIDTH - 1:0]),.Y108_out(Y108_out[2 * `WIDTH - 1:0]),.Y109_out(Y109_out[2 * `WIDTH - 1:0]),.Y110_out(Y110_out[2 * `WIDTH - 1:0]),.Y111_out(Y111_out[2 * `WIDTH - 1:0]),.Y112_out(Y112_out[2 * `WIDTH - 1:0]),
.Y113_out(Y113_out[2 * `WIDTH - 1:0]),.Y114_out(Y114_out[2 * `WIDTH - 1:0]),.Y115_out(Y115_out[2 * `WIDTH - 1:0]),.Y116_out(Y116_out[2 * `WIDTH - 1:0]),.Y117_out(Y117_out[2 * `WIDTH - 1:0]),.Y118_out(Y118_out[2 * `WIDTH - 1:0]),.Y119_out(Y119_out[2 * `WIDTH - 1:0]),.Y120_out(Y120_out[2 * `WIDTH - 1:0]),
.Y121_out(Y121_out[2 * `WIDTH - 1:0]),.Y122_out(Y122_out[2 * `WIDTH - 1:0]),.Y123_out(Y123_out[2 * `WIDTH - 1:0]),.Y124_out(Y124_out[2 * `WIDTH - 1:0]),.Y125_out(Y125_out[2 * `WIDTH - 1:0]),.Y126_out(Y126_out[2 * `WIDTH - 1:0]),.Y127_out(Y127_out[2 * `WIDTH - 1:0]),.Y128_out(Y128_out[2 * `WIDTH - 1:0]),
.Y129_out(Y129_out[2 * `WIDTH - 1:0]),.Y130_out(Y130_out[2 * `WIDTH - 1:0]),.Y131_out(Y131_out[2 * `WIDTH - 1:0]),.Y132_out(Y132_out[2 * `WIDTH - 1:0]),.Y133_out(Y133_out[2 * `WIDTH - 1:0]),.Y134_out(Y134_out[2 * `WIDTH - 1:0]),.Y135_out(Y135_out[2 * `WIDTH - 1:0]),.Y136_out(Y136_out[2 * `WIDTH - 1:0]),
.Y137_out(Y137_out[2 * `WIDTH - 1:0]),.Y138_out(Y138_out[2 * `WIDTH - 1:0]),.Y139_out(Y139_out[2 * `WIDTH - 1:0]),.Y140_out(Y140_out[2 * `WIDTH - 1:0]),.Y141_out(Y141_out[2 * `WIDTH - 1:0]),.Y142_out(Y142_out[2 * `WIDTH - 1:0]),.Y143_out(Y143_out[2 * `WIDTH - 1:0]),.Y144_out(Y144_out[2 * `WIDTH - 1:0]),
.Y145_out(Y145_out[2 * `WIDTH - 1:0]),.Y146_out(Y146_out[2 * `WIDTH - 1:0]),.Y147_out(Y147_out[2 * `WIDTH - 1:0]),.Y148_out(Y148_out[2 * `WIDTH - 1:0]),.Y149_out(Y149_out[2 * `WIDTH - 1:0]),.Y150_out(Y150_out[2 * `WIDTH - 1:0]),.Y151_out(Y151_out[2 * `WIDTH - 1:0]),.Y152_out(Y152_out[2 * `WIDTH - 1:0]),
.Y153_out(Y153_out[2 * `WIDTH - 1:0]),.Y154_out(Y154_out[2 * `WIDTH - 1:0]),.Y155_out(Y155_out[2 * `WIDTH - 1:0]),.Y156_out(Y156_out[2 * `WIDTH - 1:0]),.Y157_out(Y157_out[2 * `WIDTH - 1:0]),.Y158_out(Y158_out[2 * `WIDTH - 1:0]),.Y159_out(Y159_out[2 * `WIDTH - 1:0]),.Y160_out(Y160_out[2 * `WIDTH - 1:0]),
.Y161_out(Y161_out[2 * `WIDTH - 1:0]),.Y162_out(Y162_out[2 * `WIDTH - 1:0]),.Y163_out(Y163_out[2 * `WIDTH - 1:0]),.Y164_out(Y164_out[2 * `WIDTH - 1:0]),.Y165_out(Y165_out[2 * `WIDTH - 1:0]),.Y166_out(Y166_out[2 * `WIDTH - 1:0]),.Y167_out(Y167_out[2 * `WIDTH - 1:0]),.Y168_out(Y168_out[2 * `WIDTH - 1:0]),
.Y169_out(Y169_out[2 * `WIDTH - 1:0]),.Y170_out(Y170_out[2 * `WIDTH - 1:0]),.Y171_out(Y171_out[2 * `WIDTH - 1:0]),.Y172_out(Y172_out[2 * `WIDTH - 1:0]),.Y173_out(Y173_out[2 * `WIDTH - 1:0]),.Y174_out(Y174_out[2 * `WIDTH - 1:0]),.Y175_out(Y175_out[2 * `WIDTH - 1:0]),.Y176_out(Y176_out[2 * `WIDTH - 1:0]),
.Y177_out(Y177_out[2 * `WIDTH - 1:0]),.Y178_out(Y178_out[2 * `WIDTH - 1:0]),.Y179_out(Y179_out[2 * `WIDTH - 1:0]),.Y180_out(Y180_out[2 * `WIDTH - 1:0]),.Y181_out(Y181_out[2 * `WIDTH - 1:0]),.Y182_out(Y182_out[2 * `WIDTH - 1:0]),.Y183_out(Y183_out[2 * `WIDTH - 1:0]),.Y184_out(Y184_out[2 * `WIDTH - 1:0]),
.Y185_out(Y185_out[2 * `WIDTH - 1:0]),.Y186_out(Y186_out[2 * `WIDTH - 1:0]),.Y187_out(Y187_out[2 * `WIDTH - 1:0]),.Y188_out(Y188_out[2 * `WIDTH - 1:0]),.Y189_out(Y189_out[2 * `WIDTH - 1:0]),.Y190_out(Y190_out[2 * `WIDTH - 1:0]),.Y191_out(Y191_out[2 * `WIDTH - 1:0]),.Y192_out(Y192_out[2 * `WIDTH - 1:0]),
.Y193_out(Y193_out[2 * `WIDTH - 1:0]),.Y194_out(Y194_out[2 * `WIDTH - 1:0]),.Y195_out(Y195_out[2 * `WIDTH - 1:0]),.Y196_out(Y196_out[2 * `WIDTH - 1:0]),.Y197_out(Y197_out[2 * `WIDTH - 1:0]),.Y198_out(Y198_out[2 * `WIDTH - 1:0]),.Y199_out(Y199_out[2 * `WIDTH - 1:0]),.Y200_out(Y200_out[2 * `WIDTH - 1:0]),
.Y201_out(Y201_out[2 * `WIDTH - 1:0]),.Y202_out(Y202_out[2 * `WIDTH - 1:0]),.Y203_out(Y203_out[2 * `WIDTH - 1:0]),.Y204_out(Y204_out[2 * `WIDTH - 1:0]),.Y205_out(Y205_out[2 * `WIDTH - 1:0]),.Y206_out(Y206_out[2 * `WIDTH - 1:0]),.Y207_out(Y207_out[2 * `WIDTH - 1:0]),.Y208_out(Y208_out[2 * `WIDTH - 1:0]),
.Y209_out(Y209_out[2 * `WIDTH - 1:0]),.Y210_out(Y210_out[2 * `WIDTH - 1:0]),.Y211_out(Y211_out[2 * `WIDTH - 1:0]),.Y212_out(Y212_out[2 * `WIDTH - 1:0]),.Y213_out(Y213_out[2 * `WIDTH - 1:0]),.Y214_out(Y214_out[2 * `WIDTH - 1:0]),.Y215_out(Y215_out[2 * `WIDTH - 1:0]),.Y216_out(Y216_out[2 * `WIDTH - 1:0]),
.Y217_out(Y217_out[2 * `WIDTH - 1:0]),.Y218_out(Y218_out[2 * `WIDTH - 1:0]),.Y219_out(Y219_out[2 * `WIDTH - 1:0]),.Y220_out(Y220_out[2 * `WIDTH - 1:0]),.Y221_out(Y221_out[2 * `WIDTH - 1:0]),.Y222_out(Y222_out[2 * `WIDTH - 1:0]),.Y223_out(Y223_out[2 * `WIDTH - 1:0]),.Y224_out(Y224_out[2 * `WIDTH - 1:0]),
.Y225_out(Y225_out[2 * `WIDTH - 1:0]),.Y226_out(Y226_out[2 * `WIDTH - 1:0]),.Y227_out(Y227_out[2 * `WIDTH - 1:0]),.Y228_out(Y228_out[2 * `WIDTH - 1:0]),.Y229_out(Y229_out[2 * `WIDTH - 1:0]),.Y230_out(Y230_out[2 * `WIDTH - 1:0]),.Y231_out(Y231_out[2 * `WIDTH - 1:0]),.Y232_out(Y232_out[2 * `WIDTH - 1:0]),
.Y233_out(Y233_out[2 * `WIDTH - 1:0]),.Y234_out(Y234_out[2 * `WIDTH - 1:0]),.Y235_out(Y235_out[2 * `WIDTH - 1:0]),.Y236_out(Y236_out[2 * `WIDTH - 1:0]),.Y237_out(Y237_out[2 * `WIDTH - 1:0]),.Y238_out(Y238_out[2 * `WIDTH - 1:0]),.Y239_out(Y239_out[2 * `WIDTH - 1:0]),.Y240_out(Y240_out[2 * `WIDTH - 1:0]),
.Y241_out(Y241_out[2 * `WIDTH - 1:0]),.Y242_out(Y242_out[2 * `WIDTH - 1:0]),.Y243_out(Y243_out[2 * `WIDTH - 1:0]),.Y244_out(Y244_out[2 * `WIDTH - 1:0]),.Y245_out(Y245_out[2 * `WIDTH - 1:0]),.Y246_out(Y246_out[2 * `WIDTH - 1:0]),.Y247_out(Y247_out[2 * `WIDTH - 1:0]),.Y248_out(Y248_out[2 * `WIDTH - 1:0]),
.Y249_out(Y249_out[2 * `WIDTH - 1:0]),.Y250_out(Y250_out[2 * `WIDTH - 1:0]),.Y251_out(Y251_out[2 * `WIDTH - 1:0]),.Y252_out(Y252_out[2 * `WIDTH - 1:0]),.Y253_out(Y253_out[2 * `WIDTH - 1:0]),.Y254_out(Y254_out[2 * `WIDTH - 1:0]),.Y255_out(Y255_out[2 * `WIDTH - 1:0]),.Y256_out(Y256_out[2 * `WIDTH - 1:0]),



.I(I[`WIDTH - 1:0]),

.Initial_X_in(Initial_X[2 * `WIDTH - 1:0])
);

endmodule
