`define WIDTH 9
`define COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN 8
module sixteenbysixteen18mul (

U1_in, U2_in, U3_in, U4_in, U5_in, U6_in, U7_in, U8_in, U9_in, U10_in, U11_in, U12_in, U13_in, U14_in, U15_in, U16_in,
U17_in, U18_in, U19_in, U20_in, U21_in, U22_in, U23_in, U24_in, U25_in, U26_in, U27_in, U28_in, U29_in, U30_in, U31_in, U32_in,
U33_in, U34_in, U35_in, U36_in, U37_in, U38_in, U39_in, U40_in, U41_in, U42_in, U43_in, U44_in, U45_in, U46_in, U47_in, U48_in,
U49_in, U50_in, U51_in, U52_in, U53_in, U54_in, U55_in, U56_in, U57_in, U58_in, U59_in, U60_in, U61_in, U62_in, U63_in, U64_in,
U65_in, U66_in, U67_in, U68_in, U69_in, U70_in, U71_in, U72_in, U73_in, U74_in, U75_in, U76_in, U77_in, U78_in, U79_in, U80_in,
U81_in, U82_in, U83_in, U84_in, U85_in, U86_in, U87_in, U88_in, U89_in, U90_in, U91_in, U92_in, U93_in, U94_in, U95_in, U96_in,
U97_in, U98_in, U99_in, U100_in, U101_in, U102_in, U103_in, U104_in, U105_in, U106_in, U107_in, U108_in, U109_in, U110_in, U111_in, U112_in,
U113_in, U114_in, U115_in, U116_in, U117_in, U118_in, U119_in, U120_in, U121_in, U122_in, U123_in, U124_in, U125_in, U126_in, U127_in, U128_in,
U129_in, U130_in, U131_in, U132_in, U133_in, U134_in, U135_in, U136_in, U137_in, U138_in, U139_in, U140_in, U141_in, U142_in, U143_in, U144_in,
U145_in, U146_in, U147_in, U148_in, U149_in, U150_in, U151_in, U152_in, U153_in, U154_in, U155_in, U156_in, U157_in, U158_in, U159_in, U160_in,
U161_in, U162_in, U163_in, U164_in, U165_in, U166_in, U167_in, U168_in, U169_in, U170_in, U171_in, U172_in, U173_in, U174_in, U175_in, U176_in,
U177_in, U178_in, U179_in, U180_in, U181_in, U182_in, U183_in, U184_in, U185_in, U186_in, U187_in, U188_in, U189_in, U190_in, U191_in, U192_in,
U193_in, U194_in, U195_in, U196_in, U197_in, U198_in, U199_in, U200_in, U201_in, U202_in, U203_in, U204_in, U205_in, U206_in, U207_in, U208_in,
U209_in, U210_in, U211_in, U212_in, U213_in, U214_in, U215_in, U216_in, U217_in, U218_in, U219_in, U220_in, U221_in, U222_in, U223_in, U224_in,
U225_in, U226_in, U227_in, U228_in, U229_in, U230_in, U231_in, U232_in, U233_in, U234_in, U235_in, U236_in, U237_in, U238_in, U239_in, U240_in,
U241_in, U242_in, U243_in, U244_in, U245_in, U246_in, U247_in, U248_in, U249_in, U250_in, U251_in, U252_in, U253_in, U254_in, U255_in, U256_in,



Y1_out, Y2_out, Y3_out, Y4_out, Y5_out, Y6_out, Y7_out, Y8_out, Y9_out, Y10_out, Y11_out, Y12_out, Y13_out, Y14_out, Y15_out, Y16_out,
Y17_out, Y18_out, Y19_out, Y20_out, Y21_out, Y22_out, Y23_out, Y24_out, Y25_out, Y26_out, Y27_out, Y28_out, Y29_out, Y30_out, Y31_out, Y32_out,
Y33_out, Y34_out, Y35_out, Y36_out, Y37_out, Y38_out, Y39_out, Y40_out, Y41_out, Y42_out, Y43_out, Y44_out, Y45_out, Y46_out, Y47_out, Y48_out,
Y49_out, Y50_out, Y51_out, Y52_out, Y53_out, Y54_out, Y55_out, Y56_out, Y57_out, Y58_out, Y59_out, Y60_out, Y61_out, Y62_out, Y63_out, Y64_out,
Y65_out, Y66_out, Y67_out, Y68_out, Y69_out, Y70_out, Y71_out, Y72_out, Y73_out, Y74_out, Y75_out, Y76_out, Y77_out, Y78_out, Y79_out, Y80_out,
Y81_out, Y82_out, Y83_out, Y84_out, Y85_out, Y86_out, Y87_out, Y88_out, Y89_out, Y90_out, Y91_out, Y92_out, Y93_out, Y94_out, Y95_out, Y96_out,
Y97_out, Y98_out, Y99_out, Y100_out, Y101_out, Y102_out, Y103_out, Y104_out, Y105_out, Y106_out, Y107_out, Y108_out, Y109_out, Y110_out, Y111_out, Y112_out,
Y113_out, Y114_out, Y115_out, Y116_out, Y117_out, Y118_out, Y119_out, Y120_out, Y121_out, Y122_out, Y123_out, Y124_out, Y125_out, Y126_out, Y127_out, Y128_out,
Y129_out, Y130_out, Y131_out, Y132_out, Y133_out, Y134_out, Y135_out, Y136_out, Y137_out, Y138_out, Y139_out, Y140_out, Y141_out, Y142_out, Y143_out, Y144_out,
Y145_out, Y146_out, Y147_out, Y148_out, Y149_out, Y150_out, Y151_out, Y152_out, Y153_out, Y154_out, Y155_out, Y156_out, Y157_out, Y158_out, Y159_out, Y160_out,
Y161_out, Y162_out, Y163_out, Y164_out, Y165_out, Y166_out, Y167_out, Y168_out, Y169_out, Y170_out, Y171_out, Y172_out, Y173_out, Y174_out, Y175_out, Y176_out,
Y177_out, Y178_out, Y179_out, Y180_out, Y181_out, Y182_out, Y183_out, Y184_out, Y185_out, Y186_out, Y187_out, Y188_out, Y189_out, Y190_out, Y191_out, Y192_out,
Y193_out, Y194_out, Y195_out, Y196_out, Y197_out, Y198_out, Y199_out, Y200_out, Y201_out, Y202_out, Y203_out, Y204_out, Y205_out, Y206_out, Y207_out, Y208_out,
Y209_out, Y210_out, Y211_out, Y212_out, Y213_out, Y214_out, Y215_out, Y216_out, Y217_out, Y218_out, Y219_out, Y220_out, Y221_out, Y222_out, Y223_out, Y224_out,
Y225_out, Y226_out, Y227_out, Y228_out, Y229_out, Y230_out, Y231_out, Y232_out, Y233_out, Y234_out, Y235_out, Y236_out, Y237_out, Y238_out, Y239_out, Y240_out,
Y241_out, Y242_out, Y243_out, Y244_out, Y245_out, Y246_out, Y247_out, Y248_out, Y249_out, Y250_out, Y251_out, Y252_out, Y253_out, Y254_out, Y255_out, Y256_out,

A1, A2, A3, A4, A5, A6, A7, A8, A9,

B1, B2, B3, B4, B5, B6, B7, B8, B9,

I,

Initial_X_in,

clk
	  );
	input wire clk;
	input wire signed [`WIDTH - 1:0] I;
	input wire signed [2 * `WIDTH - 1:0] Initial_X_in;
	wire signed [2 * `WIDTH - 1:0] X_onebyoneout;
	wire signed [2 * `WIDTH - 1:0] Y_onebyoneout;
	reg signed [`WIDTH - 1:0] U1, U2, U3, U4, U5, U6, U7, U8, U9;
	reg signed [2 * `WIDTH - 1:0] Y1, Y2, Y3, Y4, Y5, Y6, Y7, Y8, Y9;
	reg [`COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN - 1:0] counter = `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b0;
	reg initial_flag = 1'b1;
	reg signed [2 * `WIDTH - 1:0] X;


	input wire signed [`WIDTH - 1:0] A1, A2, A3, A4, A5, A6, A7, A8, A9;
	input wire signed [`WIDTH - 1:0] B1, B2, B3, B4, B5, B6, B7, B8, B9;


input wire signed [`WIDTH - 1:0] U1_in, U2_in, U3_in, U4_in, U5_in, U6_in, U7_in, U8_in, U9_in, U10_in, U11_in, U12_in, U13_in, U14_in, U15_in, U16_in;
input wire signed [`WIDTH - 1:0] U17_in, U18_in, U19_in, U20_in, U21_in, U22_in, U23_in, U24_in, U25_in, U26_in, U27_in, U28_in, U29_in, U30_in, U31_in, U32_in;
input wire signed [`WIDTH - 1:0] U33_in, U34_in, U35_in, U36_in, U37_in, U38_in, U39_in, U40_in, U41_in, U42_in, U43_in, U44_in, U45_in, U46_in, U47_in, U48_in;
input wire signed [`WIDTH - 1:0] U49_in, U50_in, U51_in, U52_in, U53_in, U54_in, U55_in, U56_in, U57_in, U58_in, U59_in, U60_in, U61_in, U62_in, U63_in, U64_in;
input wire signed [`WIDTH - 1:0] U65_in, U66_in, U67_in, U68_in, U69_in, U70_in, U71_in, U72_in, U73_in, U74_in, U75_in, U76_in, U77_in, U78_in, U79_in, U80_in;
input wire signed [`WIDTH - 1:0] U81_in, U82_in, U83_in, U84_in, U85_in, U86_in, U87_in, U88_in, U89_in, U90_in, U91_in, U92_in, U93_in, U94_in, U95_in, U96_in;
input wire signed [`WIDTH - 1:0] U97_in, U98_in, U99_in, U100_in, U101_in, U102_in, U103_in, U104_in, U105_in, U106_in, U107_in, U108_in, U109_in, U110_in, U111_in, U112_in;
input wire signed [`WIDTH - 1:0] U113_in, U114_in, U115_in, U116_in, U117_in, U118_in, U119_in, U120_in, U121_in, U122_in, U123_in, U124_in, U125_in, U126_in, U127_in, U128_in;
input wire signed [`WIDTH - 1:0] U129_in, U130_in, U131_in, U132_in, U133_in, U134_in, U135_in, U136_in, U137_in, U138_in, U139_in, U140_in, U141_in, U142_in, U143_in, U144_in;
input wire signed [`WIDTH - 1:0] U145_in, U146_in, U147_in, U148_in, U149_in, U150_in, U151_in, U152_in, U153_in, U154_in, U155_in, U156_in, U157_in, U158_in, U159_in, U160_in;
input wire signed [`WIDTH - 1:0] U161_in, U162_in, U163_in, U164_in, U165_in, U166_in, U167_in, U168_in, U169_in, U170_in, U171_in, U172_in, U173_in, U174_in, U175_in, U176_in;
input wire signed [`WIDTH - 1:0] U177_in, U178_in, U179_in, U180_in, U181_in, U182_in, U183_in, U184_in, U185_in, U186_in, U187_in, U188_in, U189_in, U190_in, U191_in, U192_in;
input wire signed [`WIDTH - 1:0] U193_in, U194_in, U195_in, U196_in, U197_in, U198_in, U199_in, U200_in, U201_in, U202_in, U203_in, U204_in, U205_in, U206_in, U207_in, U208_in;
input wire signed [`WIDTH - 1:0] U209_in, U210_in, U211_in, U212_in, U213_in, U214_in, U215_in, U216_in, U217_in, U218_in, U219_in, U220_in, U221_in, U222_in, U223_in, U224_in;
input wire signed [`WIDTH - 1:0] U225_in, U226_in, U227_in, U228_in, U229_in, U230_in, U231_in, U232_in, U233_in, U234_in, U235_in, U236_in, U237_in, U238_in, U239_in, U240_in;
input wire signed [`WIDTH - 1:0] U241_in, U242_in, U243_in, U244_in, U245_in, U246_in, U247_in, U248_in, U249_in, U250_in, U251_in, U252_in, U253_in, U254_in, U255_in, U256_in;



reg signed [2 * `WIDTH - 1:0] X1_in = 0, X2_in = 0, X3_in = 0,X4_in = 0, X5_in = 0, X6_in = 0,X7_in = 0, X8_in = 0, X9_in = 0,X10_in = 0, X11_in = 0, X12_in = 0,X13_in = 0, X14_in = 0,X15_in = 0, X16_in = 0;
reg signed [2 * `WIDTH - 1:0] X17_in = 0, X18_in = 0, X19_in = 0,X20_in = 0, X21_in = 0, X22_in = 0,X23_in = 0, X24_in = 0, X25_in = 0,X26_in = 0, X27_in = 0, X28_in = 0,X29_in = 0, X30_in = 0,X31_in = 0, X32_in = 0;
reg signed [2 * `WIDTH - 1:0] X33_in = 0, X34_in = 0, X35_in = 0,X36_in = 0, X37_in = 0, X38_in = 0,X39_in = 0, X40_in = 0, X41_in = 0,X42_in = 0, X43_in = 0, X44_in = 0,X45_in = 0, X46_in = 0,X47_in = 0, X48_in = 0;
reg signed [2 * `WIDTH - 1:0] X49_in = 0, X50_in = 0, X51_in = 0,X52_in = 0, X53_in = 0, X54_in = 0,X55_in = 0, X56_in = 0, X57_in = 0,X58_in = 0, X59_in = 0, X60_in = 0,X61_in = 0, X62_in = 0,X63_in = 0, X64_in = 0;
reg signed [2 * `WIDTH - 1:0] X65_in = 0, X66_in = 0, X67_in = 0,X68_in = 0, X69_in = 0, X70_in = 0,X71_in = 0, X72_in = 0, X73_in = 0,X74_in = 0, X75_in = 0, X76_in = 0,X77_in = 0, X78_in = 0,X79_in = 0, X80_in = 0;
reg signed [2 * `WIDTH - 1:0] X81_in = 0, X82_in = 0, X83_in = 0,X84_in = 0, X85_in = 0, X86_in = 0,X87_in = 0, X88_in = 0, X89_in = 0,X90_in = 0, X91_in = 0, X92_in = 0,X93_in = 0, X94_in = 0,X95_in = 0, X96_in = 0;
reg signed [2 * `WIDTH - 1:0] X97_in = 0, X98_in = 0, X99_in = 0,X100_in = 0, X101_in = 0, X102_in = 0,X103_in = 0, X104_in = 0, X105_in = 0,X106_in = 0, X107_in = 0, X108_in = 0,X109_in = 0, X110_in = 0,X111_in = 0, X112_in = 0;
reg signed [2 * `WIDTH - 1:0] X113_in = 0, X114_in = 0, X115_in = 0,X116_in = 0, X117_in = 0, X118_in = 0,X119_in = 0, X120_in = 0, X121_in = 0,X122_in = 0, X123_in = 0, X124_in = 0,X125_in = 0, X126_in = 0,X127_in = 0, X128_in = 0;
reg signed [2 * `WIDTH - 1:0] X129_in = 0, X130_in = 0, X131_in = 0,X132_in = 0, X133_in = 0, X134_in = 0,X135_in = 0, X136_in = 0, X137_in = 0,X138_in = 0, X139_in = 0, X140_in = 0,X141_in = 0, X142_in = 0,X143_in = 0, X144_in = 0;
reg signed [2 * `WIDTH - 1:0] X145_in = 0, X146_in = 0, X147_in = 0,X148_in = 0, X149_in = 0, X150_in = 0,X151_in = 0, X152_in = 0, X153_in = 0,X154_in = 0, X155_in = 0, X156_in = 0,X157_in = 0, X158_in = 0,X159_in = 0, X160_in = 0;
reg signed [2 * `WIDTH - 1:0] X161_in = 0, X162_in = 0, X163_in = 0,X164_in = 0, X165_in = 0, X166_in = 0,X167_in = 0, X168_in = 0, X169_in = 0,X170_in = 0, X171_in = 0, X172_in = 0,X173_in = 0, X174_in = 0,X175_in = 0, X176_in = 0;
reg signed [2 * `WIDTH - 1:0] X177_in = 0, X178_in = 0, X179_in = 0,X180_in = 0, X181_in = 0, X182_in = 0,X183_in = 0, X184_in = 0, X185_in = 0,X186_in = 0, X187_in = 0, X188_in = 0,X189_in = 0, X190_in = 0,X191_in = 0, X192_in = 0;
reg signed [2 * `WIDTH - 1:0] X193_in = 0, X194_in = 0, X195_in = 0,X196_in = 0, X197_in = 0, X198_in = 0,X199_in = 0, X200_in = 0, X201_in = 0,X202_in = 0, X203_in = 0, X204_in = 0,X205_in = 0, X206_in = 0,X207_in = 0, X208_in = 0;
reg signed [2 * `WIDTH - 1:0] X209_in = 0, X210_in = 0, X211_in = 0,X212_in = 0, X213_in = 0, X214_in = 0,X215_in = 0, X216_in = 0, X217_in = 0,X218_in = 0, X219_in = 0, X220_in = 0,X221_in = 0, X222_in = 0,X223_in = 0, X224_in = 0;
reg signed [2 * `WIDTH - 1:0] X225_in = 0, X226_in = 0, X227_in = 0,X228_in = 0, X229_in = 0, X230_in = 0,X231_in = 0, X232_in = 0, X233_in = 0,X234_in = 0, X235_in = 0, X236_in = 0,X237_in = 0, X238_in = 0,X239_in = 0, X240_in = 0;
reg signed [2 * `WIDTH - 1:0] X241_in = 0, X242_in = 0, X243_in = 0,X244_in = 0, X245_in = 0, X246_in = 0,X247_in = 0, X248_in = 0, X249_in = 0,X250_in = 0, X251_in = 0, X252_in = 0,X253_in = 0, X254_in = 0,X255_in = 0, X256_in = 0;



reg signed [2 * `WIDTH - 1:0] X1_next = 0, X2_next = 0, X3_next = 0,X4_next = 0, X5_next = 0, X6_next = 0,X7_next = 0, X8_next = 0, X9_next = 0,X10_next = 0, X11_next = 0, X12_next = 0,X13_next = 0, X14_next = 0,X15_next = 0, X16_next = 0;
reg signed [2 * `WIDTH - 1:0] X17_next = 0, X18_next = 0, X19_next = 0,X20_next = 0, X21_next = 0, X22_next = 0,X23_next = 0, X24_next = 0, X25_next = 0,X26_next = 0, X27_next = 0, X28_next = 0,X29_next = 0, X30_next = 0,X31_next = 0, X32_next = 0;
reg signed [2 * `WIDTH - 1:0] X33_next = 0, X34_next = 0, X35_next = 0,X36_next = 0, X37_next = 0, X38_next = 0,X39_next = 0, X40_next = 0, X41_next = 0,X42_next = 0, X43_next = 0, X44_next = 0,X45_next = 0, X46_next = 0,X47_next = 0, X48_next = 0;
reg signed [2 * `WIDTH - 1:0] X49_next = 0, X50_next = 0, X51_next = 0,X52_next = 0, X53_next = 0, X54_next = 0,X55_next = 0, X56_next = 0, X57_next = 0,X58_next = 0, X59_next = 0, X60_next = 0,X61_next = 0, X62_next = 0,X63_next = 0, X64_next = 0;
reg signed [2 * `WIDTH - 1:0] X65_next = 0, X66_next = 0, X67_next = 0,X68_next = 0, X69_next = 0, X70_next = 0,X71_next = 0, X72_next = 0, X73_next = 0,X74_next = 0, X75_next = 0, X76_next = 0,X77_next = 0, X78_next = 0,X79_next = 0, X80_next = 0;
reg signed [2 * `WIDTH - 1:0] X81_next = 0, X82_next = 0, X83_next = 0,X84_next = 0, X85_next = 0, X86_next = 0,X87_next = 0, X88_next = 0, X89_next = 0,X90_next = 0, X91_next = 0, X92_next = 0,X93_next = 0, X94_next = 0,X95_next = 0, X96_next = 0;
reg signed [2 * `WIDTH - 1:0] X97_next = 0, X98_next = 0, X99_next = 0,X100_next = 0, X101_next = 0, X102_next = 0,X103_next = 0, X104_next = 0, X105_next = 0,X106_next = 0, X107_next = 0, X108_next = 0,X109_next = 0, X110_next = 0,X111_next = 0, X112_next = 0;
reg signed [2 * `WIDTH - 1:0] X113_next = 0, X114_next = 0, X115_next = 0,X116_next = 0, X117_next = 0, X118_next = 0,X119_next = 0, X120_next = 0, X121_next = 0,X122_next = 0, X123_next = 0, X124_next = 0,X125_next = 0, X126_next = 0,X127_next = 0, X128_next = 0;
reg signed [2 * `WIDTH - 1:0] X129_next = 0, X130_next = 0, X131_next = 0,X132_next = 0, X133_next = 0, X134_next = 0,X135_next = 0, X136_next = 0, X137_next = 0,X138_next = 0, X139_next = 0, X140_next = 0,X141_next = 0, X142_next = 0,X143_next = 0, X144_next = 0;
reg signed [2 * `WIDTH - 1:0] X145_next = 0, X146_next = 0, X147_next = 0,X148_next = 0, X149_next = 0, X150_next = 0,X151_next = 0, X152_next = 0, X153_next = 0,X154_next = 0, X155_next = 0, X156_next = 0,X157_next = 0, X158_next = 0,X159_next = 0, X160_next = 0;
reg signed [2 * `WIDTH - 1:0] X161_next = 0, X162_next = 0, X163_next = 0,X164_next = 0, X165_next = 0, X166_next = 0,X167_next = 0, X168_next = 0, X169_next = 0,X170_next = 0, X171_next = 0, X172_next = 0,X173_next = 0, X174_next = 0,X175_next = 0, X176_next = 0;
reg signed [2 * `WIDTH - 1:0] X177_next = 0, X178_next = 0, X179_next = 0,X180_next = 0, X181_next = 0, X182_next = 0,X183_next = 0, X184_next = 0, X185_next = 0,X186_next = 0, X187_next = 0, X188_next = 0,X189_next = 0, X190_next = 0,X191_next = 0, X192_next = 0;
reg signed [2 * `WIDTH - 1:0] X193_next = 0, X194_next = 0, X195_next = 0,X196_next = 0, X197_next = 0, X198_next = 0,X199_next = 0, X200_next = 0, X201_next = 0,X202_next = 0, X203_next = 0, X204_next = 0,X205_next = 0, X206_next = 0,X207_next = 0, X208_next = 0;
reg signed [2 * `WIDTH - 1:0] X209_next = 0, X210_next = 0, X211_next = 0,X212_next = 0, X213_next = 0, X214_next = 0,X215_next = 0, X216_next = 0, X217_next = 0,X218_next = 0, X219_next = 0, X220_next = 0,X221_next = 0, X222_next = 0,X223_next = 0, X224_next = 0;
reg signed [2 * `WIDTH - 1:0] X225_next = 0, X226_next = 0, X227_next = 0,X228_next = 0, X229_next = 0, X230_next = 0,X231_next = 0, X232_next = 0, X233_next = 0,X234_next = 0, X235_next = 0, X236_next = 0,X237_next = 0, X238_next = 0,X239_next = 0, X240_next = 0;
reg signed [2 * `WIDTH - 1:0] X241_next = 0, X242_next = 0, X243_next = 0,X244_next = 0, X245_next = 0, X246_next = 0,X247_next = 0, X248_next = 0, X249_next = 0,X250_next = 0, X251_next = 0, X252_next = 0,X253_next = 0, X254_next = 0,X255_next = 0, X256_next = 0;



reg signed [2 * `WIDTH - 1:0] Y1_in = 0, Y2_in = 0, Y3_in = 0,Y4_in = 0, Y5_in = 0, Y6_in = 0,Y7_in = 0, Y8_in = 0, Y9_in = 0,Y10_in = 0, Y11_in = 0, Y12_in = 0,Y13_in = 0, Y14_in = 0,Y15_in = 0, Y16_in = 0;
reg signed [2 * `WIDTH - 1:0] Y17_in = 0, Y18_in = 0, Y19_in = 0,Y20_in = 0, Y21_in = 0, Y22_in = 0,Y23_in = 0, Y24_in = 0, Y25_in = 0,Y26_in = 0, Y27_in = 0, Y28_in = 0,Y29_in = 0, Y30_in = 0,Y31_in = 0, Y32_in = 0;
reg signed [2 * `WIDTH - 1:0] Y33_in = 0, Y34_in = 0, Y35_in = 0,Y36_in = 0, Y37_in = 0, Y38_in = 0,Y39_in = 0, Y40_in = 0, Y41_in = 0,Y42_in = 0, Y43_in = 0, Y44_in = 0,Y45_in = 0, Y46_in = 0,Y47_in = 0, Y48_in = 0;
reg signed [2 * `WIDTH - 1:0] Y49_in = 0, Y50_in = 0, Y51_in = 0,Y52_in = 0, Y53_in = 0, Y54_in = 0,Y55_in = 0, Y56_in = 0, Y57_in = 0,Y58_in = 0, Y59_in = 0, Y60_in = 0,Y61_in = 0, Y62_in = 0,Y63_in = 0, Y64_in = 0;
reg signed [2 * `WIDTH - 1:0] Y65_in = 0, Y66_in = 0, Y67_in = 0,Y68_in = 0, Y69_in = 0, Y70_in = 0,Y71_in = 0, Y72_in = 0, Y73_in = 0,Y74_in = 0, Y75_in = 0, Y76_in = 0,Y77_in = 0, Y78_in = 0,Y79_in = 0, Y80_in = 0;
reg signed [2 * `WIDTH - 1:0] Y81_in = 0, Y82_in = 0, Y83_in = 0,Y84_in = 0, Y85_in = 0, Y86_in = 0,Y87_in = 0, Y88_in = 0, Y89_in = 0,Y90_in = 0, Y91_in = 0, Y92_in = 0,Y93_in = 0, Y94_in = 0,Y95_in = 0, Y96_in = 0;
reg signed [2 * `WIDTH - 1:0] Y97_in = 0, Y98_in = 0, Y99_in = 0,Y100_in = 0, Y101_in = 0, Y102_in = 0,Y103_in = 0, Y104_in = 0, Y105_in = 0,Y106_in = 0, Y107_in = 0, Y108_in = 0,Y109_in = 0, Y110_in = 0,Y111_in = 0, Y112_in = 0;
reg signed [2 * `WIDTH - 1:0] Y113_in = 0, Y114_in = 0, Y115_in = 0,Y116_in = 0, Y117_in = 0, Y118_in = 0,Y119_in = 0, Y120_in = 0, Y121_in = 0,Y122_in = 0, Y123_in = 0, Y124_in = 0,Y125_in = 0, Y126_in = 0,Y127_in = 0, Y128_in = 0;
reg signed [2 * `WIDTH - 1:0] Y129_in = 0, Y130_in = 0, Y131_in = 0,Y132_in = 0, Y133_in = 0, Y134_in = 0,Y135_in = 0, Y136_in = 0, Y137_in = 0,Y138_in = 0, Y139_in = 0, Y140_in = 0,Y141_in = 0, Y142_in = 0,Y143_in = 0, Y144_in = 0;
reg signed [2 * `WIDTH - 1:0] Y145_in = 0, Y146_in = 0, Y147_in = 0,Y148_in = 0, Y149_in = 0, Y150_in = 0,Y151_in = 0, Y152_in = 0, Y153_in = 0,Y154_in = 0, Y155_in = 0, Y156_in = 0,Y157_in = 0, Y158_in = 0,Y159_in = 0, Y160_in = 0;
reg signed [2 * `WIDTH - 1:0] Y161_in = 0, Y162_in = 0, Y163_in = 0,Y164_in = 0, Y165_in = 0, Y166_in = 0,Y167_in = 0, Y168_in = 0, Y169_in = 0,Y170_in = 0, Y171_in = 0, Y172_in = 0,Y173_in = 0, Y174_in = 0,Y175_in = 0, Y176_in = 0;
reg signed [2 * `WIDTH - 1:0] Y177_in = 0, Y178_in = 0, Y179_in = 0,Y180_in = 0, Y181_in = 0, Y182_in = 0,Y183_in = 0, Y184_in = 0, Y185_in = 0,Y186_in = 0, Y187_in = 0, Y188_in = 0,Y189_in = 0, Y190_in = 0,Y191_in = 0, Y192_in = 0;
reg signed [2 * `WIDTH - 1:0] Y193_in = 0, Y194_in = 0, Y195_in = 0,Y196_in = 0, Y197_in = 0, Y198_in = 0,Y199_in = 0, Y200_in = 0, Y201_in = 0,Y202_in = 0, Y203_in = 0, Y204_in = 0,Y205_in = 0, Y206_in = 0,Y207_in = 0, Y208_in = 0;
reg signed [2 * `WIDTH - 1:0] Y209_in = 0, Y210_in = 0, Y211_in = 0,Y212_in = 0, Y213_in = 0, Y214_in = 0,Y215_in = 0, Y216_in = 0, Y217_in = 0,Y218_in = 0, Y219_in = 0, Y220_in = 0,Y221_in = 0, Y222_in = 0,Y223_in = 0, Y224_in = 0;
reg signed [2 * `WIDTH - 1:0] Y225_in = 0, Y226_in = 0, Y227_in = 0,Y228_in = 0, Y229_in = 0, Y230_in = 0,Y231_in = 0, Y232_in = 0, Y233_in = 0,Y234_in = 0, Y235_in = 0, Y236_in = 0,Y237_in = 0, Y238_in = 0,Y239_in = 0, Y240_in = 0;
reg signed [2 * `WIDTH - 1:0] Y241_in = 0, Y242_in = 0, Y243_in = 0,Y244_in = 0, Y245_in = 0, Y246_in = 0,Y247_in = 0, Y248_in = 0, Y249_in = 0,Y250_in = 0, Y251_in = 0, Y252_in = 0,Y253_in = 0, Y254_in = 0,Y255_in = 0, Y256_in = 0;



reg signed [2 * `WIDTH - 1:0] Y1_next = 0, Y2_next = 0, Y3_next = 0,Y4_next = 0, Y5_next = 0, Y6_next = 0,Y7_next = 0, Y8_next = 0, Y9_next = 0,Y10_next = 0, Y11_next = 0, Y12_next = 0,Y13_next = 0, Y14_next = 0,Y15_next = 0, Y16_next = 0;
reg signed [2 * `WIDTH - 1:0] Y17_next = 0, Y18_next = 0, Y19_next = 0,Y20_next = 0, Y21_next = 0, Y22_next = 0,Y23_next = 0, Y24_next = 0, Y25_next = 0,Y26_next = 0, Y27_next = 0, Y28_next = 0,Y29_next = 0, Y30_next = 0,Y31_next = 0, Y32_next = 0;
reg signed [2 * `WIDTH - 1:0] Y33_next = 0, Y34_next = 0, Y35_next = 0,Y36_next = 0, Y37_next = 0, Y38_next = 0,Y39_next = 0, Y40_next = 0, Y41_next = 0,Y42_next = 0, Y43_next = 0, Y44_next = 0,Y45_next = 0, Y46_next = 0,Y47_next = 0, Y48_next = 0;
reg signed [2 * `WIDTH - 1:0] Y49_next = 0, Y50_next = 0, Y51_next = 0,Y52_next = 0, Y53_next = 0, Y54_next = 0,Y55_next = 0, Y56_next = 0, Y57_next = 0,Y58_next = 0, Y59_next = 0, Y60_next = 0,Y61_next = 0, Y62_next = 0,Y63_next = 0, Y64_next = 0;
reg signed [2 * `WIDTH - 1:0] Y65_next = 0, Y66_next = 0, Y67_next = 0,Y68_next = 0, Y69_next = 0, Y70_next = 0,Y71_next = 0, Y72_next = 0, Y73_next = 0,Y74_next = 0, Y75_next = 0, Y76_next = 0,Y77_next = 0, Y78_next = 0,Y79_next = 0, Y80_next = 0;
reg signed [2 * `WIDTH - 1:0] Y81_next = 0, Y82_next = 0, Y83_next = 0,Y84_next = 0, Y85_next = 0, Y86_next = 0,Y87_next = 0, Y88_next = 0, Y89_next = 0,Y90_next = 0, Y91_next = 0, Y92_next = 0,Y93_next = 0, Y94_next = 0,Y95_next = 0, Y96_next = 0;
reg signed [2 * `WIDTH - 1:0] Y97_next = 0, Y98_next = 0, Y99_next = 0,Y100_next = 0, Y101_next = 0, Y102_next = 0,Y103_next = 0, Y104_next = 0, Y105_next = 0,Y106_next = 0, Y107_next = 0, Y108_next = 0,Y109_next = 0, Y110_next = 0,Y111_next = 0, Y112_next = 0;
reg signed [2 * `WIDTH - 1:0] Y113_next = 0, Y114_next = 0, Y115_next = 0,Y116_next = 0, Y117_next = 0, Y118_next = 0,Y119_next = 0, Y120_next = 0, Y121_next = 0,Y122_next = 0, Y123_next = 0, Y124_next = 0,Y125_next = 0, Y126_next = 0,Y127_next = 0, Y128_next = 0;
reg signed [2 * `WIDTH - 1:0] Y129_next = 0, Y130_next = 0, Y131_next = 0,Y132_next = 0, Y133_next = 0, Y134_next = 0,Y135_next = 0, Y136_next = 0, Y137_next = 0,Y138_next = 0, Y139_next = 0, Y140_next = 0,Y141_next = 0, Y142_next = 0,Y143_next = 0, Y144_next = 0;
reg signed [2 * `WIDTH - 1:0] Y145_next = 0, Y146_next = 0, Y147_next = 0,Y148_next = 0, Y149_next = 0, Y150_next = 0,Y151_next = 0, Y152_next = 0, Y153_next = 0,Y154_next = 0, Y155_next = 0, Y156_next = 0,Y157_next = 0, Y158_next = 0,Y159_next = 0, Y160_next = 0;
reg signed [2 * `WIDTH - 1:0] Y161_next = 0, Y162_next = 0, Y163_next = 0,Y164_next = 0, Y165_next = 0, Y166_next = 0,Y167_next = 0, Y168_next = 0, Y169_next = 0,Y170_next = 0, Y171_next = 0, Y172_next = 0,Y173_next = 0, Y174_next = 0,Y175_next = 0, Y176_next = 0;
reg signed [2 * `WIDTH - 1:0] Y177_next = 0, Y178_next = 0, Y179_next = 0,Y180_next = 0, Y181_next = 0, Y182_next = 0,Y183_next = 0, Y184_next = 0, Y185_next = 0,Y186_next = 0, Y187_next = 0, Y188_next = 0,Y189_next = 0, Y190_next = 0,Y191_next = 0, Y192_next = 0;
reg signed [2 * `WIDTH - 1:0] Y193_next = 0, Y194_next = 0, Y195_next = 0,Y196_next = 0, Y197_next = 0, Y198_next = 0,Y199_next = 0, Y200_next = 0, Y201_next = 0,Y202_next = 0, Y203_next = 0, Y204_next = 0,Y205_next = 0, Y206_next = 0,Y207_next = 0, Y208_next = 0;
reg signed [2 * `WIDTH - 1:0] Y209_next = 0, Y210_next = 0, Y211_next = 0,Y212_next = 0, Y213_next = 0, Y214_next = 0,Y215_next = 0, Y216_next = 0, Y217_next = 0,Y218_next = 0, Y219_next = 0, Y220_next = 0,Y221_next = 0, Y222_next = 0,Y223_next = 0, Y224_next = 0;
reg signed [2 * `WIDTH - 1:0] Y225_next = 0, Y226_next = 0, Y227_next = 0,Y228_next = 0, Y229_next = 0, Y230_next = 0,Y231_next = 0, Y232_next = 0, Y233_next = 0,Y234_next = 0, Y235_next = 0, Y236_next = 0,Y237_next = 0, Y238_next = 0,Y239_next = 0, Y240_next = 0;
reg signed [2 * `WIDTH - 1:0] Y241_next = 0, Y242_next = 0, Y243_next = 0,Y244_next = 0, Y245_next = 0, Y246_next = 0,Y247_next = 0, Y248_next = 0, Y249_next = 0,Y250_next = 0, Y251_next = 0, Y252_next = 0,Y253_next = 0, Y254_next = 0,Y255_next = 0, Y256_next = 0;



output wire signed [2 * `WIDTH - 1:0] Y1_out, Y2_out, Y3_out, Y4_out, Y5_out, Y6_out, Y7_out, Y8_out, Y9_out, Y10_out, Y11_out, Y12_out, Y13_out, Y14_out, Y15_out, Y16_out;
output wire signed [2 * `WIDTH - 1:0] Y17_out, Y18_out, Y19_out, Y20_out, Y21_out, Y22_out, Y23_out, Y24_out, Y25_out, Y26_out, Y27_out, Y28_out, Y29_out, Y30_out, Y31_out, Y32_out;
output wire signed [2 * `WIDTH - 1:0] Y33_out, Y34_out, Y35_out, Y36_out, Y37_out, Y38_out, Y39_out, Y40_out, Y41_out, Y42_out, Y43_out, Y44_out, Y45_out, Y46_out, Y47_out, Y48_out;
output wire signed [2 * `WIDTH - 1:0] Y49_out, Y50_out, Y51_out, Y52_out, Y53_out, Y54_out, Y55_out, Y56_out, Y57_out, Y58_out, Y59_out, Y60_out, Y61_out, Y62_out, Y63_out, Y64_out;
output wire signed [2 * `WIDTH - 1:0] Y65_out, Y66_out, Y67_out, Y68_out, Y69_out, Y70_out, Y71_out, Y72_out, Y73_out, Y74_out, Y75_out, Y76_out, Y77_out, Y78_out, Y79_out, Y80_out;
output wire signed [2 * `WIDTH - 1:0] Y81_out, Y82_out, Y83_out, Y84_out, Y85_out, Y86_out, Y87_out, Y88_out, Y89_out, Y90_out, Y91_out, Y92_out, Y93_out, Y94_out, Y95_out, Y96_out;
output wire signed [2 * `WIDTH - 1:0] Y97_out, Y98_out, Y99_out, Y100_out, Y101_out, Y102_out, Y103_out, Y104_out, Y105_out, Y106_out, Y107_out, Y108_out, Y109_out, Y110_out, Y111_out, Y112_out;
output wire signed [2 * `WIDTH - 1:0] Y113_out, Y114_out, Y115_out, Y116_out, Y117_out, Y118_out, Y119_out, Y120_out, Y121_out, Y122_out, Y123_out, Y124_out, Y125_out, Y126_out, Y127_out, Y128_out;
output wire signed [2 * `WIDTH - 1:0] Y129_out, Y130_out, Y131_out, Y132_out, Y133_out, Y134_out, Y135_out, Y136_out, Y137_out, Y138_out, Y139_out, Y140_out, Y141_out, Y142_out, Y143_out, Y144_out;
output wire signed [2 * `WIDTH - 1:0] Y145_out, Y146_out, Y147_out, Y148_out, Y149_out, Y150_out, Y151_out, Y152_out, Y153_out, Y154_out, Y155_out, Y156_out, Y157_out, Y158_out, Y159_out, Y160_out;
output wire signed [2 * `WIDTH - 1:0] Y161_out, Y162_out, Y163_out, Y164_out, Y165_out, Y166_out, Y167_out, Y168_out, Y169_out, Y170_out, Y171_out, Y172_out, Y173_out, Y174_out, Y175_out, Y176_out;
output wire signed [2 * `WIDTH - 1:0] Y177_out, Y178_out, Y179_out, Y180_out, Y181_out, Y182_out, Y183_out, Y184_out, Y185_out, Y186_out, Y187_out, Y188_out, Y189_out, Y190_out, Y191_out, Y192_out;
output wire signed [2 * `WIDTH - 1:0] Y193_out, Y194_out, Y195_out, Y196_out, Y197_out, Y198_out, Y199_out, Y200_out, Y201_out, Y202_out, Y203_out, Y204_out, Y205_out, Y206_out, Y207_out, Y208_out;
output wire signed [2 * `WIDTH - 1:0] Y209_out, Y210_out, Y211_out, Y212_out, Y213_out, Y214_out, Y215_out, Y216_out, Y217_out, Y218_out, Y219_out, Y220_out, Y221_out, Y222_out, Y223_out, Y224_out;
output wire signed [2 * `WIDTH - 1:0] Y225_out, Y226_out, Y227_out, Y228_out, Y229_out, Y230_out, Y231_out, Y232_out, Y233_out, Y234_out, Y235_out, Y236_out, Y237_out, Y238_out, Y239_out, Y240_out;
output wire signed [2 * `WIDTH - 1:0] Y241_out, Y242_out, Y243_out, Y244_out, Y245_out, Y246_out, Y247_out, Y248_out, Y249_out, Y250_out, Y251_out, Y252_out, Y253_out, Y254_out, Y255_out, Y256_out;



assign Y1_out = Y1_next;assign Y2_out = Y2_next;assign Y3_out = Y3_next;assign Y4_out = Y4_next;assign Y5_out = Y5_next;assign Y6_out = Y6_next;assign Y7_out = Y7_next;assign Y8_out = Y8_next;
assign Y9_out = Y9_next;assign Y10_out = Y10_next;assign Y11_out = Y11_next;assign Y12_out = Y12_next;assign Y13_out = Y13_next;assign Y14_out = Y14_next;assign Y15_out = Y15_next;assign Y16_out = Y16_next;
assign Y17_out = Y17_next;assign Y18_out = Y18_next;assign Y19_out = Y19_next;assign Y20_out = Y20_next;assign Y21_out = Y21_next;assign Y22_out = Y22_next;assign Y23_out = Y23_next;assign Y24_out = Y24_next;
assign Y25_out = Y25_next;assign Y26_out = Y26_next;assign Y27_out = Y27_next;assign Y28_out = Y28_next;assign Y29_out = Y29_next;assign Y30_out = Y30_next;assign Y31_out = Y31_next;assign Y32_out = Y32_next;
assign Y33_out = Y33_next;assign Y34_out = Y34_next;assign Y35_out = Y35_next;assign Y36_out = Y36_next;assign Y37_out = Y37_next;assign Y38_out = Y38_next;assign Y39_out = Y39_next;assign Y40_out = Y40_next;
assign Y41_out = Y41_next;assign Y42_out = Y42_next;assign Y43_out = Y43_next;assign Y44_out = Y44_next;assign Y45_out = Y45_next;assign Y46_out = Y46_next;assign Y47_out = Y47_next;assign Y48_out = Y48_next;
assign Y49_out = Y49_next;assign Y50_out = Y50_next;assign Y51_out = Y51_next;assign Y52_out = Y52_next;assign Y53_out = Y53_next;assign Y54_out = Y54_next;assign Y55_out = Y55_next;assign Y56_out = Y56_next;
assign Y57_out = Y57_next;assign Y58_out = Y58_next;assign Y59_out = Y59_next;assign Y60_out = Y60_next;assign Y61_out = Y61_next;assign Y62_out = Y62_next;assign Y63_out = Y63_next;assign Y64_out = Y64_next;
assign Y65_out = Y65_next;assign Y66_out = Y66_next;assign Y67_out = Y67_next;assign Y68_out = Y68_next;assign Y69_out = Y69_next;assign Y70_out = Y70_next;assign Y71_out = Y71_next;assign Y72_out = Y72_next;
assign Y73_out = Y73_next;assign Y74_out = Y74_next;assign Y75_out = Y75_next;assign Y76_out = Y76_next;assign Y77_out = Y77_next;assign Y78_out = Y78_next;assign Y79_out = Y79_next;assign Y80_out = Y80_next;
assign Y81_out = Y81_next;assign Y82_out = Y82_next;assign Y83_out = Y83_next;assign Y84_out = Y84_next;assign Y85_out = Y85_next;assign Y86_out = Y86_next;assign Y87_out = Y87_next;assign Y88_out = Y88_next;
assign Y89_out = Y89_next;assign Y90_out = Y90_next;assign Y91_out = Y91_next;assign Y92_out = Y92_next;assign Y93_out = Y93_next;assign Y94_out = Y94_next;assign Y95_out = Y95_next;assign Y96_out = Y96_next;
assign Y97_out = Y97_next;assign Y98_out = Y98_next;assign Y99_out = Y99_next;assign Y100_out = Y100_next;assign Y101_out = Y101_next;assign Y102_out = Y102_next;assign Y103_out = Y103_next;assign Y104_out = Y104_next;
assign Y105_out = Y105_next;assign Y106_out = Y106_next;assign Y107_out = Y107_next;assign Y108_out = Y108_next;assign Y109_out = Y109_next;assign Y110_out = Y110_next;assign Y111_out = Y111_next;assign Y112_out = Y112_next;
assign Y113_out = Y113_next;assign Y114_out = Y114_next;assign Y115_out = Y115_next;assign Y116_out = Y116_next;assign Y117_out = Y117_next;assign Y118_out = Y118_next;assign Y119_out = Y119_next;assign Y120_out = Y120_next;
assign Y121_out = Y121_next;assign Y122_out = Y122_next;assign Y123_out = Y123_next;assign Y124_out = Y124_next;assign Y125_out = Y125_next;assign Y126_out = Y126_next;assign Y127_out = Y127_next;assign Y128_out = Y128_next;
assign Y129_out = Y129_next;assign Y130_out = Y130_next;assign Y131_out = Y131_next;assign Y132_out = Y132_next;assign Y133_out = Y133_next;assign Y134_out = Y134_next;assign Y135_out = Y135_next;assign Y136_out = Y136_next;
assign Y137_out = Y137_next;assign Y138_out = Y138_next;assign Y139_out = Y139_next;assign Y140_out = Y140_next;assign Y141_out = Y141_next;assign Y142_out = Y142_next;assign Y143_out = Y143_next;assign Y144_out = Y144_next;
assign Y145_out = Y145_next;assign Y146_out = Y146_next;assign Y147_out = Y147_next;assign Y148_out = Y148_next;assign Y149_out = Y149_next;assign Y150_out = Y150_next;assign Y151_out = Y151_next;assign Y152_out = Y152_next;
assign Y153_out = Y153_next;assign Y154_out = Y154_next;assign Y155_out = Y155_next;assign Y156_out = Y156_next;assign Y157_out = Y157_next;assign Y158_out = Y158_next;assign Y159_out = Y159_next;assign Y160_out = Y160_next;
assign Y161_out = Y161_next;assign Y162_out = Y162_next;assign Y163_out = Y163_next;assign Y164_out = Y164_next;assign Y165_out = Y165_next;assign Y166_out = Y166_next;assign Y167_out = Y167_next;assign Y168_out = Y168_next;
assign Y169_out = Y169_next;assign Y170_out = Y170_next;assign Y171_out = Y171_next;assign Y172_out = Y172_next;assign Y173_out = Y173_next;assign Y174_out = Y174_next;assign Y175_out = Y175_next;assign Y176_out = Y176_next;
assign Y177_out = Y177_next;assign Y178_out = Y178_next;assign Y179_out = Y179_next;assign Y180_out = Y180_next;assign Y181_out = Y181_next;assign Y182_out = Y182_next;assign Y183_out = Y183_next;assign Y184_out = Y184_next;
assign Y185_out = Y185_next;assign Y186_out = Y186_next;assign Y187_out = Y187_next;assign Y188_out = Y188_next;assign Y189_out = Y189_next;assign Y190_out = Y190_next;assign Y191_out = Y191_next;assign Y192_out = Y192_next;
assign Y193_out = Y193_next;assign Y194_out = Y194_next;assign Y195_out = Y195_next;assign Y196_out = Y196_next;assign Y197_out = Y197_next;assign Y198_out = Y198_next;assign Y199_out = Y199_next;assign Y200_out = Y200_next;
assign Y201_out = Y201_next;assign Y202_out = Y202_next;assign Y203_out = Y203_next;assign Y204_out = Y204_next;assign Y205_out = Y205_next;assign Y206_out = Y206_next;assign Y207_out = Y207_next;assign Y208_out = Y208_next;
assign Y209_out = Y209_next;assign Y210_out = Y210_next;assign Y211_out = Y211_next;assign Y212_out = Y212_next;assign Y213_out = Y213_next;assign Y214_out = Y214_next;assign Y215_out = Y215_next;assign Y216_out = Y216_next;
assign Y217_out = Y217_next;assign Y218_out = Y218_next;assign Y219_out = Y219_next;assign Y220_out = Y220_next;assign Y221_out = Y221_next;assign Y222_out = Y222_next;assign Y223_out = Y223_next;assign Y224_out = Y224_next;
assign Y225_out = Y225_next;assign Y226_out = Y226_next;assign Y227_out = Y227_next;assign Y228_out = Y228_next;assign Y229_out = Y229_next;assign Y230_out = Y230_next;assign Y231_out = Y231_next;assign Y232_out = Y232_next;
assign Y233_out = Y233_next;assign Y234_out = Y234_next;assign Y235_out = Y235_next;assign Y236_out = Y236_next;assign Y237_out = Y237_next;assign Y238_out = Y238_next;assign Y239_out = Y239_next;assign Y240_out = Y240_next;
assign Y241_out = Y241_next;assign Y242_out = Y242_next;assign Y243_out = Y243_next;assign Y244_out = Y244_next;assign Y245_out = Y245_next;assign Y246_out = Y246_next;assign Y247_out = Y247_next;assign Y248_out = Y248_next;
assign Y249_out = Y249_next;assign Y250_out = Y250_next;assign Y251_out = Y251_next;assign Y252_out = Y252_next;assign Y253_out = Y253_next;assign Y254_out = Y254_next;assign Y255_out = Y255_next;assign Y256_out = Y256_next;





always  @ (posedge clk)
begin
  if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b0) begin // 1

	if (initial_flag == 1'b0) begin

		Y256_next <= Y_onebyoneout;
		X256_next <= X_onebyoneout;

Y1_in = Y1_next;Y2_in = Y2_next;Y3_in = Y3_next;Y4_in = Y4_next;Y5_in = Y5_next;Y6_in = Y6_next;Y7_in = Y7_next;Y8_in = Y8_next;
Y9_in = Y9_next;Y10_in = Y10_next;Y11_in = Y11_next;Y12_in = Y12_next;Y13_in = Y13_next;Y14_in = Y14_next;Y15_in = Y15_next;Y16_in = Y16_next;
Y17_in = Y17_next;Y18_in = Y18_next;Y19_in = Y19_next;Y20_in = Y20_next;Y21_in = Y21_next;Y22_in = Y22_next;Y23_in = Y23_next;Y24_in = Y24_next;
Y25_in = Y25_next;Y26_in = Y26_next;Y27_in = Y27_next;Y28_in = Y28_next;Y29_in = Y29_next;Y30_in = Y30_next;Y31_in = Y31_next;Y32_in = Y32_next;
Y33_in = Y33_next;Y34_in = Y34_next;Y35_in = Y35_next;Y36_in = Y36_next;Y37_in = Y37_next;Y38_in = Y38_next;Y39_in = Y39_next;Y40_in = Y40_next;
Y41_in = Y41_next;Y42_in = Y42_next;Y43_in = Y43_next;Y44_in = Y44_next;Y45_in = Y45_next;Y46_in = Y46_next;Y47_in = Y47_next;Y48_in = Y48_next;
Y49_in = Y49_next;Y50_in = Y50_next;Y51_in = Y51_next;Y52_in = Y52_next;Y53_in = Y53_next;Y54_in = Y54_next;Y55_in = Y55_next;Y56_in = Y56_next;
Y57_in = Y57_next;Y58_in = Y58_next;Y59_in = Y59_next;Y60_in = Y60_next;Y61_in = Y61_next;Y62_in = Y62_next;Y63_in = Y63_next;Y64_in = Y64_next;
Y65_in = Y65_next;Y66_in = Y66_next;Y67_in = Y67_next;Y68_in = Y68_next;Y69_in = Y69_next;Y70_in = Y70_next;Y71_in = Y71_next;Y72_in = Y72_next;
Y73_in = Y73_next;Y74_in = Y74_next;Y75_in = Y75_next;Y76_in = Y76_next;Y77_in = Y77_next;Y78_in = Y78_next;Y79_in = Y79_next;Y80_in = Y80_next;
Y81_in = Y81_next;Y82_in = Y82_next;Y83_in = Y83_next;Y84_in = Y84_next;Y85_in = Y85_next;Y86_in = Y86_next;Y87_in = Y87_next;Y88_in = Y88_next;
Y89_in = Y89_next;Y90_in = Y90_next;Y91_in = Y91_next;Y92_in = Y92_next;Y93_in = Y93_next;Y94_in = Y94_next;Y95_in = Y95_next;Y96_in = Y96_next;
Y97_in = Y97_next;Y98_in = Y98_next;Y99_in = Y99_next;Y100_in = Y100_next;Y101_in = Y101_next;Y102_in = Y102_next;Y103_in = Y103_next;Y104_in = Y104_next;
Y105_in = Y105_next;Y106_in = Y106_next;Y107_in = Y107_next;Y108_in = Y108_next;Y109_in = Y109_next;Y110_in = Y110_next;Y111_in = Y111_next;Y112_in = Y112_next;
Y113_in = Y113_next;Y114_in = Y114_next;Y115_in = Y115_next;Y116_in = Y116_next;Y117_in = Y117_next;Y118_in = Y118_next;Y119_in = Y119_next;Y120_in = Y120_next;
Y121_in = Y121_next;Y122_in = Y122_next;Y123_in = Y123_next;Y124_in = Y124_next;Y125_in = Y125_next;Y126_in = Y126_next;Y127_in = Y127_next;Y128_in = Y128_next;
Y129_in = Y129_next;Y130_in = Y130_next;Y131_in = Y131_next;Y132_in = Y132_next;Y133_in = Y133_next;Y134_in = Y134_next;Y135_in = Y135_next;Y136_in = Y136_next;
Y137_in = Y137_next;Y138_in = Y138_next;Y139_in = Y139_next;Y140_in = Y140_next;Y141_in = Y141_next;Y142_in = Y142_next;Y143_in = Y143_next;Y144_in = Y144_next;
Y145_in = Y145_next;Y146_in = Y146_next;Y147_in = Y147_next;Y148_in = Y148_next;Y149_in = Y149_next;Y150_in = Y150_next;Y151_in = Y151_next;Y152_in = Y152_next;
Y153_in = Y153_next;Y154_in = Y154_next;Y155_in = Y155_next;Y156_in = Y156_next;Y157_in = Y157_next;Y158_in = Y158_next;Y159_in = Y159_next;Y160_in = Y160_next;
Y161_in = Y161_next;Y162_in = Y162_next;Y163_in = Y163_next;Y164_in = Y164_next;Y165_in = Y165_next;Y166_in = Y166_next;Y167_in = Y167_next;Y168_in = Y168_next;
Y169_in = Y169_next;Y170_in = Y170_next;Y171_in = Y171_next;Y172_in = Y172_next;Y173_in = Y173_next;Y174_in = Y174_next;Y175_in = Y175_next;Y176_in = Y176_next;
Y177_in = Y177_next;Y178_in = Y178_next;Y179_in = Y179_next;Y180_in = Y180_next;Y181_in = Y181_next;Y182_in = Y182_next;Y183_in = Y183_next;Y184_in = Y184_next;
Y185_in = Y185_next;Y186_in = Y186_next;Y187_in = Y187_next;Y188_in = Y188_next;Y189_in = Y189_next;Y190_in = Y190_next;Y191_in = Y191_next;Y192_in = Y192_next;
Y193_in = Y193_next;Y194_in = Y194_next;Y195_in = Y195_next;Y196_in = Y196_next;Y197_in = Y197_next;Y198_in = Y198_next;Y199_in = Y199_next;Y200_in = Y200_next;
Y201_in = Y201_next;Y202_in = Y202_next;Y203_in = Y203_next;Y204_in = Y204_next;Y205_in = Y205_next;Y206_in = Y206_next;Y207_in = Y207_next;Y208_in = Y208_next;
Y209_in = Y209_next;Y210_in = Y210_next;Y211_in = Y211_next;Y212_in = Y212_next;Y213_in = Y213_next;Y214_in = Y214_next;Y215_in = Y215_next;Y216_in = Y216_next;
Y217_in = Y217_next;Y218_in = Y218_next;Y219_in = Y219_next;Y220_in = Y220_next;Y221_in = Y221_next;Y222_in = Y222_next;Y223_in = Y223_next;Y224_in = Y224_next;
Y225_in = Y225_next;Y226_in = Y226_next;Y227_in = Y227_next;Y228_in = Y228_next;Y229_in = Y229_next;Y230_in = Y230_next;Y231_in = Y231_next;Y232_in = Y232_next;
Y233_in = Y233_next;Y234_in = Y234_next;Y235_in = Y235_next;Y236_in = Y236_next;Y237_in = Y237_next;Y238_in = Y238_next;Y239_in = Y239_next;Y240_in = Y240_next;
Y241_in = Y241_next;Y242_in = Y242_next;Y243_in = Y243_next;Y244_in = Y244_next;Y245_in = Y245_next;Y246_in = Y246_next;Y247_in = Y247_next;Y248_in = Y248_next;
Y249_in = Y249_next;Y250_in = Y250_next;Y251_in = Y251_next;Y252_in = Y252_next;Y253_in = Y253_next;Y254_in = Y254_next;Y255_in = Y255_next;Y256_in = Y256_next;

X1_in = X1_next;X2_in = X2_next;X3_in = X3_next;X4_in = X4_next;X5_in = X5_next;X6_in = X6_next;X7_in = X7_next;X8_in = X8_next;
X9_in = X9_next;X10_in = X10_next;X11_in = X11_next;X12_in = X12_next;X13_in = X13_next;X14_in = X14_next;X15_in = X15_next;X16_in = X16_next;
X17_in = X17_next;X18_in = X18_next;X19_in = X19_next;X20_in = X20_next;X21_in = X21_next;X22_in = X22_next;X23_in = X23_next;X24_in = X24_next;
X25_in = X25_next;X26_in = X26_next;X27_in = X27_next;X28_in = X28_next;X29_in = X29_next;X30_in = X30_next;X31_in = X31_next;X32_in = X32_next;
X33_in = X33_next;X34_in = X34_next;X35_in = X35_next;X36_in = X36_next;X37_in = X37_next;X38_in = X38_next;X39_in = X39_next;X40_in = X40_next;
X41_in = X41_next;X42_in = X42_next;X43_in = X43_next;X44_in = X44_next;X45_in = X45_next;X46_in = X46_next;X47_in = X47_next;X48_in = X48_next;
X49_in = X49_next;X50_in = X50_next;X51_in = X51_next;X52_in = X52_next;X53_in = X53_next;X54_in = X54_next;X55_in = X55_next;X56_in = X56_next;
X57_in = X57_next;X58_in = X58_next;X59_in = X59_next;X60_in = X60_next;X61_in = X61_next;X62_in = X62_next;X63_in = X63_next;X64_in = X64_next;
X65_in = X65_next;X66_in = X66_next;X67_in = X67_next;X68_in = X68_next;X69_in = X69_next;X70_in = X70_next;X71_in = X71_next;X72_in = X72_next;
X73_in = X73_next;X74_in = X74_next;X75_in = X75_next;X76_in = X76_next;X77_in = X77_next;X78_in = X78_next;X79_in = X79_next;X80_in = X80_next;
X81_in = X81_next;X82_in = X82_next;X83_in = X83_next;X84_in = X84_next;X85_in = X85_next;X86_in = X86_next;X87_in = X87_next;X88_in = X88_next;
X89_in = X89_next;X90_in = X90_next;X91_in = X91_next;X92_in = X92_next;X93_in = X93_next;X94_in = X94_next;X95_in = X95_next;X96_in = X96_next;
X97_in = X97_next;X98_in = X98_next;X99_in = X99_next;X100_in = X100_next;X101_in = X101_next;X102_in = X102_next;X103_in = X103_next;X104_in = X104_next;
X105_in = X105_next;X106_in = X106_next;X107_in = X107_next;X108_in = X108_next;X109_in = X109_next;X110_in = X110_next;X111_in = X111_next;X112_in = X112_next;
X113_in = X113_next;X114_in = X114_next;X115_in = X115_next;X116_in = X116_next;X117_in = X117_next;X118_in = X118_next;X119_in = X119_next;X120_in = X120_next;
X121_in = X121_next;X122_in = X122_next;X123_in = X123_next;X124_in = X124_next;X125_in = X125_next;X126_in = X126_next;X127_in = X127_next;X128_in = X128_next;
X129_in = X129_next;X130_in = X130_next;X131_in = X131_next;X132_in = X132_next;X133_in = X133_next;X134_in = X134_next;X135_in = X135_next;X136_in = X136_next;
X137_in = X137_next;X138_in = X138_next;X139_in = X139_next;X140_in = X140_next;X141_in = X141_next;X142_in = X142_next;X143_in = X143_next;X144_in = X144_next;
X145_in = X145_next;X146_in = X146_next;X147_in = X147_next;X148_in = X148_next;X149_in = X149_next;X150_in = X150_next;X151_in = X151_next;X152_in = X152_next;
X153_in = X153_next;X154_in = X154_next;X155_in = X155_next;X156_in = X156_next;X157_in = X157_next;X158_in = X158_next;X159_in = X159_next;X160_in = X160_next;
X161_in = X161_next;X162_in = X162_next;X163_in = X163_next;X164_in = X164_next;X165_in = X165_next;X166_in = X166_next;X167_in = X167_next;X168_in = X168_next;
X169_in = X169_next;X170_in = X170_next;X171_in = X171_next;X172_in = X172_next;X173_in = X173_next;X174_in = X174_next;X175_in = X175_next;X176_in = X176_next;
X177_in = X177_next;X178_in = X178_next;X179_in = X179_next;X180_in = X180_next;X181_in = X181_next;X182_in = X182_next;X183_in = X183_next;X184_in = X184_next;
X185_in = X185_next;X186_in = X186_next;X187_in = X187_next;X188_in = X188_next;X189_in = X189_next;X190_in = X190_next;X191_in = X191_next;X192_in = X192_next;
X193_in = X193_next;X194_in = X194_next;X195_in = X195_next;X196_in = X196_next;X197_in = X197_next;X198_in = X198_next;X199_in = X199_next;X200_in = X200_next;
X201_in = X201_next;X202_in = X202_next;X203_in = X203_next;X204_in = X204_next;X205_in = X205_next;X206_in = X206_next;X207_in = X207_next;X208_in = X208_next;
X209_in = X209_next;X210_in = X210_next;X211_in = X211_next;X212_in = X212_next;X213_in = X213_next;X214_in = X214_next;X215_in = X215_next;X216_in = X216_next;
X217_in = X217_next;X218_in = X218_next;X219_in = X219_next;X220_in = X220_next;X221_in = X221_next;X222_in = X222_next;X223_in = X223_next;X224_in = X224_next;
X225_in = X225_next;X226_in = X226_next;X227_in = X227_next;X228_in = X228_next;X229_in = X229_next;X230_in = X230_next;X231_in = X231_next;X232_in = X232_next;
X233_in = X233_next;X234_in = X234_next;X235_in = X235_next;X236_in = X236_next;X237_in = X237_next;X238_in = X238_next;X239_in = X239_next;X240_in = X240_next;
X241_in = X241_next;X242_in = X242_next;X243_in = X243_next;X244_in = X244_next;X245_in = X245_next;X246_in = X246_next;X247_in = X247_next;X248_in = X248_next;
X249_in = X249_next;X250_in = X250_next;X251_in = X251_next;X252_in = X252_next;X253_in = X253_next;X254_in = X254_next;X255_in = X255_next;X256_in = X256_next;

	end else begin

X1_in = Initial_X_in;X2_in = Initial_X_in;X3_in = Initial_X_in;X4_in = Initial_X_in;X5_in = Initial_X_in;X6_in = Initial_X_in;X7_in = Initial_X_in; X8_in = Initial_X_in;
X9_in = Initial_X_in;X10_in = Initial_X_in;X11_in = Initial_X_in;X12_in = Initial_X_in;X13_in = Initial_X_in;X14_in = Initial_X_in;X15_in = Initial_X_in; X16_in = Initial_X_in;
X17_in = Initial_X_in;X18_in = Initial_X_in;X19_in = Initial_X_in;X20_in = Initial_X_in;X21_in = Initial_X_in;X22_in = Initial_X_in;X23_in = Initial_X_in; X24_in = Initial_X_in;
X25_in = Initial_X_in;X26_in = Initial_X_in;X27_in = Initial_X_in;X28_in = Initial_X_in;X29_in = Initial_X_in;X30_in = Initial_X_in;X31_in = Initial_X_in; X32_in = Initial_X_in;
X33_in = Initial_X_in;X34_in = Initial_X_in;X35_in = Initial_X_in;X36_in = Initial_X_in;X37_in = Initial_X_in;X38_in = Initial_X_in;X39_in = Initial_X_in; X40_in = Initial_X_in;
X41_in = Initial_X_in;X42_in = Initial_X_in;X43_in = Initial_X_in;X44_in = Initial_X_in;X45_in = Initial_X_in;X46_in = Initial_X_in;X47_in = Initial_X_in; X48_in = Initial_X_in;
X49_in = Initial_X_in;X50_in = Initial_X_in;X51_in = Initial_X_in;X52_in = Initial_X_in;X53_in = Initial_X_in;X54_in = Initial_X_in;X55_in = Initial_X_in; X56_in = Initial_X_in;
X57_in = Initial_X_in;X58_in = Initial_X_in;X59_in = Initial_X_in;X60_in = Initial_X_in;X61_in = Initial_X_in;X62_in = Initial_X_in;X63_in = Initial_X_in; X64_in = Initial_X_in;
X65_in = Initial_X_in;X66_in = Initial_X_in;X67_in = Initial_X_in;X68_in = Initial_X_in;X69_in = Initial_X_in;X70_in = Initial_X_in;X71_in = Initial_X_in; X72_in = Initial_X_in;
X73_in = Initial_X_in;X74_in = Initial_X_in;X75_in = Initial_X_in;X76_in = Initial_X_in;X77_in = Initial_X_in;X78_in = Initial_X_in;X79_in = Initial_X_in; X80_in = Initial_X_in;
X81_in = Initial_X_in;X82_in = Initial_X_in;X83_in = Initial_X_in;X84_in = Initial_X_in;X85_in = Initial_X_in;X86_in = Initial_X_in;X87_in = Initial_X_in; X88_in = Initial_X_in;
X89_in = Initial_X_in;X90_in = Initial_X_in;X91_in = Initial_X_in;X92_in = Initial_X_in;X93_in = Initial_X_in;X94_in = Initial_X_in;X95_in = Initial_X_in; X96_in = Initial_X_in;
X97_in = Initial_X_in;X98_in = Initial_X_in;X99_in = Initial_X_in;X100_in = Initial_X_in;X101_in = Initial_X_in;X102_in = Initial_X_in;X103_in = Initial_X_in; X104_in = Initial_X_in;
X105_in = Initial_X_in;X106_in = Initial_X_in;X107_in = Initial_X_in;X108_in = Initial_X_in;X109_in = Initial_X_in;X110_in = Initial_X_in;X111_in = Initial_X_in; X112_in = Initial_X_in;
X113_in = Initial_X_in;X114_in = Initial_X_in;X115_in = Initial_X_in;X116_in = Initial_X_in;X117_in = Initial_X_in;X118_in = Initial_X_in;X119_in = Initial_X_in; X120_in = Initial_X_in;
X121_in = Initial_X_in;X122_in = Initial_X_in;X123_in = Initial_X_in;X124_in = Initial_X_in;X125_in = Initial_X_in;X126_in = Initial_X_in;X127_in = Initial_X_in; X128_in = Initial_X_in;
X129_in = Initial_X_in;X130_in = Initial_X_in;X131_in = Initial_X_in;X132_in = Initial_X_in;X133_in = Initial_X_in;X134_in = Initial_X_in;X135_in = Initial_X_in; X136_in = Initial_X_in;
X137_in = Initial_X_in;X138_in = Initial_X_in;X139_in = Initial_X_in;X140_in = Initial_X_in;X141_in = Initial_X_in;X142_in = Initial_X_in;X143_in = Initial_X_in; X144_in = Initial_X_in;
X145_in = Initial_X_in;X146_in = Initial_X_in;X147_in = Initial_X_in;X148_in = Initial_X_in;X149_in = Initial_X_in;X150_in = Initial_X_in;X151_in = Initial_X_in; X152_in = Initial_X_in;
X153_in = Initial_X_in;X154_in = Initial_X_in;X155_in = Initial_X_in;X156_in = Initial_X_in;X157_in = Initial_X_in;X158_in = Initial_X_in;X159_in = Initial_X_in; X160_in = Initial_X_in;
X161_in = Initial_X_in;X162_in = Initial_X_in;X163_in = Initial_X_in;X164_in = Initial_X_in;X165_in = Initial_X_in;X166_in = Initial_X_in;X167_in = Initial_X_in; X168_in = Initial_X_in;
X169_in = Initial_X_in;X170_in = Initial_X_in;X171_in = Initial_X_in;X172_in = Initial_X_in;X173_in = Initial_X_in;X174_in = Initial_X_in;X175_in = Initial_X_in; X176_in = Initial_X_in;
X177_in = Initial_X_in;X178_in = Initial_X_in;X179_in = Initial_X_in;X180_in = Initial_X_in;X181_in = Initial_X_in;X182_in = Initial_X_in;X183_in = Initial_X_in; X184_in = Initial_X_in;
X185_in = Initial_X_in;X186_in = Initial_X_in;X187_in = Initial_X_in;X188_in = Initial_X_in;X189_in = Initial_X_in;X190_in = Initial_X_in;X191_in = Initial_X_in; X192_in = Initial_X_in;
X193_in = Initial_X_in;X194_in = Initial_X_in;X195_in = Initial_X_in;X196_in = Initial_X_in;X197_in = Initial_X_in;X198_in = Initial_X_in;X199_in = Initial_X_in; X200_in = Initial_X_in;
X201_in = Initial_X_in;X202_in = Initial_X_in;X203_in = Initial_X_in;X204_in = Initial_X_in;X205_in = Initial_X_in;X206_in = Initial_X_in;X207_in = Initial_X_in; X208_in = Initial_X_in;
X209_in = Initial_X_in;X210_in = Initial_X_in;X211_in = Initial_X_in;X212_in = Initial_X_in;X213_in = Initial_X_in;X214_in = Initial_X_in;X215_in = Initial_X_in; X216_in = Initial_X_in;
X217_in = Initial_X_in;X218_in = Initial_X_in;X219_in = Initial_X_in;X220_in = Initial_X_in;X221_in = Initial_X_in;X222_in = Initial_X_in;X223_in = Initial_X_in; X224_in = Initial_X_in;
X225_in = Initial_X_in;X226_in = Initial_X_in;X227_in = Initial_X_in;X228_in = Initial_X_in;X229_in = Initial_X_in;X230_in = Initial_X_in;X231_in = Initial_X_in; X232_in = Initial_X_in;
X233_in = Initial_X_in;X234_in = Initial_X_in;X235_in = Initial_X_in;X236_in = Initial_X_in;X237_in = Initial_X_in;X238_in = Initial_X_in;X239_in = Initial_X_in; X240_in = Initial_X_in;
X241_in = Initial_X_in;X242_in = Initial_X_in;X243_in = Initial_X_in;X244_in = Initial_X_in;X245_in = Initial_X_in;X246_in = Initial_X_in;X247_in = Initial_X_in; X248_in = Initial_X_in;
X249_in = Initial_X_in;X250_in = Initial_X_in;X251_in = Initial_X_in;X252_in = Initial_X_in;X253_in = Initial_X_in;X254_in = Initial_X_in;X255_in = Initial_X_in; X256_in = Initial_X_in;

		initial_flag = 1'b0;
	end

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= `WIDTH'b0;
    U5 <= U1_in;
    U6 <= U2_in;
    U7 <= `WIDTH'b0;
    U8 <= U17_in;
    U9 <= U18_in;

    X <= X1_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y1_in;
    Y6 <= Y2_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y17_in;
    Y9 <= Y18_in;

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1) begin // 2

    Y1_next <= Y_onebyoneout;
    X1_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U1_in;
    U5 <= U2_in;
    U6 <= U3_in;
    U7 <= U17_in;
    U8 <= U18_in;
    U9 <= U19_in;

    X <= X2_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y1_in;
    Y5 <= Y2_in;
    Y6 <= Y3_in;
    Y7 <= Y17_in;
    Y8 <= Y18_in;
    Y9 <= Y19_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10) begin // 3

    Y2_next <= Y_onebyoneout;
    X2_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U2_in;
    U5 <= U3_in;
    U6 <= U4_in;
    U7 <= U18_in;
    U8 <= U19_in;
    U9 <= U20_in;

    X <= X3_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y2_in;
    Y5 <= Y3_in;
    Y6 <= Y4_in;
    Y7 <= Y18_in;
    Y8 <= Y19_in;
    Y9 <= Y20_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11) begin // 4

    Y3_next <= Y_onebyoneout;
    X3_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U3_in;
    U5 <= U4_in;
    U6 <= U5_in;
    U7 <= U19_in;
    U8 <= U20_in;
    U9 <= U21_in;

    X <= X4_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y3_in;
    Y5 <= Y4_in;
    Y6 <= Y5_in;
    Y7 <= Y19_in;
    Y8 <= Y20_in;
    Y9 <= Y21_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b100) begin // 5

    Y4_next <= Y_onebyoneout;
    X4_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U4_in;
    U5 <= U5_in;
    U6 <= U6_in;
    U7 <= U20_in;
    U8 <= U21_in;
    U9 <= U22_in;

    X <= X5_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y4_in;
    Y5 <= Y5_in;
    Y6 <= Y6_in;
    Y7 <= Y20_in;
    Y8 <= Y21_in;
    Y9 <= Y22_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b101) begin // 6

    Y5_next <= Y_onebyoneout;
    X5_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U5_in;
    U5 <= U6_in;
    U6 <= U7_in;
    U7 <= U21_in;
    U8 <= U22_in;
    U9 <= U23_in;

    X <= X6_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y5_in;
    Y5 <= Y6_in;
    Y6 <= Y7_in;
    Y7 <= Y21_in;
    Y8 <= Y22_in;
    Y9 <= Y23_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b110) begin // 7

    Y6_next <= Y_onebyoneout;
    X6_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U6_in;
    U5 <= U7_in;
    U6 <= U8_in;
    U7 <= U22_in;
    U8 <= U23_in;
    U9 <= U24_in;

    X <= X7_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y6_in;
    Y5 <= Y7_in;
    Y6 <= Y8_in;
    Y7 <= Y22_in;
    Y8 <= Y23_in;
    Y9 <= Y24_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b111) begin // 8

    Y7_next <= Y_onebyoneout;
    X7_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U7_in;
    U5 <= U8_in;
    U6 <= U9_in;
    U7 <= U23_in;
    U8 <= U24_in;
    U9 <= U25_in;

    X <= X8_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y7_in;
    Y5 <= Y8_in;
    Y6 <= Y9_in;
    Y7 <= Y23_in;
    Y8 <= Y24_in;
    Y9 <= Y25_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1000) begin // 9

    Y8_next <= Y_onebyoneout;
    X8_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U8_in;
    U5 <= U9_in;
    U6 <= U10_in;
    U7 <= U24_in;
    U8 <= U25_in;
    U9 <= U26_in;

    X <= X9_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y8_in;
    Y5 <= Y9_in;
    Y6 <= Y10_in;
    Y7 <= Y24_in;
    Y8 <= Y25_in;
    Y9 <= Y26_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1001) begin // 10

    Y9_next <= Y_onebyoneout;
    X9_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U9_in;
    U5 <= U10_in;
    U6 <= U11_in;
    U7 <= U25_in;
    U8 <= U26_in;
    U9 <= U27_in;

    X <= X10_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y9_in;
    Y5 <= Y10_in;
    Y6 <= Y11_in;
    Y7 <= Y25_in;
    Y8 <= Y26_in;
    Y9 <= Y27_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1010) begin // 11

    Y10_next <= Y_onebyoneout;
    X10_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U10_in;
    U5 <= U11_in;
    U6 <= U12_in;
    U7 <= U26_in;
    U8 <= U27_in;
    U9 <= U28_in;

    X <= X11_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y10_in;
    Y5 <= Y11_in;
    Y6 <= Y12_in;
    Y7 <= Y26_in;
    Y8 <= Y27_in;
    Y9 <= Y28_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1011) begin // 12

    Y11_next <= Y_onebyoneout;
    X11_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U11_in;
    U5 <= U12_in;
    U6 <= U13_in;
    U7 <= U27_in;
    U8 <= U28_in;
    U9 <= U29_in;

    X <= X12_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y11_in;
    Y5 <= Y12_in;
    Y6 <= Y13_in;
    Y7 <= Y27_in;
    Y8 <= Y28_in;
    Y9 <= Y29_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1100) begin // 13

    Y12_next <= Y_onebyoneout;
    X12_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U12_in;
    U5 <= U13_in;
    U6 <= U14_in;
    U7 <= U28_in;
    U8 <= U29_in;
    U9 <= U30_in;

    X <= X13_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y12_in;
    Y5 <= Y13_in;
    Y6 <= Y14_in;
    Y7 <= Y28_in;
    Y8 <= Y29_in;
    Y9 <= Y30_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1101) begin // 14

    Y13_next <= Y_onebyoneout;
    X13_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U13_in;
    U5 <= U14_in;
    U6 <= U15_in;
    U7 <= U29_in;
    U8 <= U30_in;
    U9 <= U31_in;

    X <= X14_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y13_in;
    Y5 <= Y14_in;
    Y6 <= Y15_in;
    Y7 <= Y29_in;
    Y8 <= Y30_in;
    Y9 <= Y31_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1110) begin // 15

    Y14_next <= Y_onebyoneout;
    X14_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U14_in;
    U5 <= U15_in;
    U6 <= U16_in;
    U7 <= U30_in;
    U8 <= U31_in;
    U9 <= U32_in;

    X <= X15_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y14_in;
    Y5 <= Y15_in;
    Y6 <= Y16_in;
    Y7 <= Y30_in;
    Y8 <= Y31_in;
    Y9 <= Y32_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1111) begin // 16

    Y15_next <= Y_onebyoneout;
    X15_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= `WIDTH'b0;
    U3 <= `WIDTH'b0;
    U4 <= U15_in;
    U5 <= U16_in;
    U6 <= `WIDTH'b0;
    U7 <= U31_in;
    U8 <= U32_in;
    U9 <= `WIDTH'b0;

    X <= X16_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= {(2 * `WIDTH){1'b0}};
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y15_in;
    Y5 <= Y16_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y31_in;
    Y8 <= Y32_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10000) begin // 17

    Y16_next <= Y_onebyoneout;
    X16_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U1_in;
    U3 <= U2_in;
    U4 <= `WIDTH'b0;
    U5 <= U17_in;
    U6 <= U18_in;
    U7 <= `WIDTH'b0;
    U8 <= U33_in;
    U9 <= U34_in;

    X <= X17_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y1_in;
    Y3 <= Y2_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y17_in;
    Y6 <= Y18_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y33_in;
    Y9 <= Y34_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10001) begin // 18

    Y17_next <= Y_onebyoneout;
    X17_next <= X_onebyoneout;

    U1 <= U1_in;
    U2 <= U2_in;
    U3 <= U3_in;
    U4 <= U17_in;
    U5 <= U18_in;
    U6 <= U19_in;
    U7 <= U33_in;
    U8 <= U34_in;
    U9 <= U35_in;

    X <= X18_in;

    Y1 <= Y1_in;
    Y2 <= Y2_in;
    Y3 <= Y3_in;
    Y4 <= Y17_in;
    Y5 <= Y18_in;
    Y6 <= Y19_in;
    Y7 <= Y33_in;
    Y8 <= Y34_in;
    Y9 <= Y35_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10010) begin // 19

    Y18_next <= Y_onebyoneout;
    X18_next <= X_onebyoneout;

    U1 <= U2_in;
    U2 <= U3_in;
    U3 <= U4_in;
    U4 <= U18_in;
    U5 <= U19_in;
    U6 <= U20_in;
    U7 <= U34_in;
    U8 <= U35_in;
    U9 <= U36_in;

    X <= X19_in;

    Y1 <= Y2_in;
    Y2 <= Y3_in;
    Y3 <= Y4_in;
    Y4 <= Y18_in;
    Y5 <= Y19_in;
    Y6 <= Y20_in;
    Y7 <= Y34_in;
    Y8 <= Y35_in;
    Y9 <= Y36_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10011) begin // 20

    Y19_next <= Y_onebyoneout;
    X19_next <= X_onebyoneout;

    U1 <= U3_in;
    U2 <= U4_in;
    U3 <= U5_in;
    U4 <= U19_in;
    U5 <= U20_in;
    U6 <= U21_in;
    U7 <= U35_in;
    U8 <= U36_in;
    U9 <= U37_in;

    X <= X20_in;

    Y1 <= Y3_in;
    Y2 <= Y4_in;
    Y3 <= Y5_in;
    Y4 <= Y19_in;
    Y5 <= Y20_in;
    Y6 <= Y21_in;
    Y7 <= Y35_in;
    Y8 <= Y36_in;
    Y9 <= Y37_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10100) begin // 21

    Y20_next <= Y_onebyoneout;
    X20_next <= X_onebyoneout;

    U1 <= U4_in;
    U2 <= U5_in;
    U3 <= U6_in;
    U4 <= U20_in;
    U5 <= U21_in;
    U6 <= U22_in;
    U7 <= U36_in;
    U8 <= U37_in;
    U9 <= U38_in;

    X <= X21_in;

    Y1 <= Y4_in;
    Y2 <= Y5_in;
    Y3 <= Y6_in;
    Y4 <= Y20_in;
    Y5 <= Y21_in;
    Y6 <= Y22_in;
    Y7 <= Y36_in;
    Y8 <= Y37_in;
    Y9 <= Y38_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10101) begin // 22

    Y21_next <= Y_onebyoneout;
    X21_next <= X_onebyoneout;

    U1 <= U5_in;
    U2 <= U6_in;
    U3 <= U7_in;
    U4 <= U21_in;
    U5 <= U22_in;
    U6 <= U23_in;
    U7 <= U37_in;
    U8 <= U38_in;
    U9 <= U39_in;

    X <= X22_in;

    Y1 <= Y5_in;
    Y2 <= Y6_in;
    Y3 <= Y7_in;
    Y4 <= Y21_in;
    Y5 <= Y22_in;
    Y6 <= Y23_in;
    Y7 <= Y37_in;
    Y8 <= Y38_in;
    Y9 <= Y39_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10110) begin // 23

    Y22_next <= Y_onebyoneout;
    X22_next <= X_onebyoneout;

    U1 <= U6_in;
    U2 <= U7_in;
    U3 <= U8_in;
    U4 <= U22_in;
    U5 <= U23_in;
    U6 <= U24_in;
    U7 <= U38_in;
    U8 <= U39_in;
    U9 <= U40_in;

    X <= X23_in;

    Y1 <= Y6_in;
    Y2 <= Y7_in;
    Y3 <= Y8_in;
    Y4 <= Y22_in;
    Y5 <= Y23_in;
    Y6 <= Y24_in;
    Y7 <= Y38_in;
    Y8 <= Y39_in;
    Y9 <= Y40_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10111) begin // 24

    Y23_next <= Y_onebyoneout;
    X23_next <= X_onebyoneout;

    U1 <= U7_in;
    U2 <= U8_in;
    U3 <= U9_in;
    U4 <= U23_in;
    U5 <= U24_in;
    U6 <= U25_in;
    U7 <= U39_in;
    U8 <= U40_in;
    U9 <= U41_in;

    X <= X24_in;

    Y1 <= Y7_in;
    Y2 <= Y8_in;
    Y3 <= Y9_in;
    Y4 <= Y23_in;
    Y5 <= Y24_in;
    Y6 <= Y25_in;
    Y7 <= Y39_in;
    Y8 <= Y40_in;
    Y9 <= Y41_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11000) begin // 25

    Y24_next <= Y_onebyoneout;
    X24_next <= X_onebyoneout;

    U1 <= U8_in;
    U2 <= U9_in;
    U3 <= U10_in;
    U4 <= U24_in;
    U5 <= U25_in;
    U6 <= U26_in;
    U7 <= U40_in;
    U8 <= U41_in;
    U9 <= U42_in;

    X <= X25_in;

    Y1 <= Y8_in;
    Y2 <= Y9_in;
    Y3 <= Y10_in;
    Y4 <= Y24_in;
    Y5 <= Y25_in;
    Y6 <= Y26_in;
    Y7 <= Y40_in;
    Y8 <= Y41_in;
    Y9 <= Y42_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11001) begin // 26

    Y25_next <= Y_onebyoneout;
    X25_next <= X_onebyoneout;

    U1 <= U9_in;
    U2 <= U10_in;
    U3 <= U11_in;
    U4 <= U25_in;
    U5 <= U26_in;
    U6 <= U27_in;
    U7 <= U41_in;
    U8 <= U42_in;
    U9 <= U43_in;

    X <= X26_in;

    Y1 <= Y9_in;
    Y2 <= Y10_in;
    Y3 <= Y11_in;
    Y4 <= Y25_in;
    Y5 <= Y26_in;
    Y6 <= Y27_in;
    Y7 <= Y41_in;
    Y8 <= Y42_in;
    Y9 <= Y43_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11010) begin // 27

    Y26_next <= Y_onebyoneout;
    X26_next <= X_onebyoneout;

    U1 <= U10_in;
    U2 <= U11_in;
    U3 <= U12_in;
    U4 <= U26_in;
    U5 <= U27_in;
    U6 <= U28_in;
    U7 <= U42_in;
    U8 <= U43_in;
    U9 <= U44_in;

    X <= X27_in;

    Y1 <= Y10_in;
    Y2 <= Y11_in;
    Y3 <= Y12_in;
    Y4 <= Y26_in;
    Y5 <= Y27_in;
    Y6 <= Y28_in;
    Y7 <= Y42_in;
    Y8 <= Y43_in;
    Y9 <= Y44_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11011) begin // 28

    Y27_next <= Y_onebyoneout;
    X27_next <= X_onebyoneout;

    U1 <= U11_in;
    U2 <= U12_in;
    U3 <= U13_in;
    U4 <= U27_in;
    U5 <= U28_in;
    U6 <= U29_in;
    U7 <= U43_in;
    U8 <= U44_in;
    U9 <= U45_in;

    X <= X28_in;

    Y1 <= Y11_in;
    Y2 <= Y12_in;
    Y3 <= Y13_in;
    Y4 <= Y27_in;
    Y5 <= Y28_in;
    Y6 <= Y29_in;
    Y7 <= Y43_in;
    Y8 <= Y44_in;
    Y9 <= Y45_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11100) begin // 29

    Y28_next <= Y_onebyoneout;
    X28_next <= X_onebyoneout;

    U1 <= U12_in;
    U2 <= U13_in;
    U3 <= U14_in;
    U4 <= U28_in;
    U5 <= U29_in;
    U6 <= U30_in;
    U7 <= U44_in;
    U8 <= U45_in;
    U9 <= U46_in;

    X <= X29_in;

    Y1 <= Y12_in;
    Y2 <= Y13_in;
    Y3 <= Y14_in;
    Y4 <= Y28_in;
    Y5 <= Y29_in;
    Y6 <= Y30_in;
    Y7 <= Y44_in;
    Y8 <= Y45_in;
    Y9 <= Y46_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11101) begin // 30

    Y29_next <= Y_onebyoneout;
    X29_next <= X_onebyoneout;

    U1 <= U13_in;
    U2 <= U14_in;
    U3 <= U15_in;
    U4 <= U29_in;
    U5 <= U30_in;
    U6 <= U31_in;
    U7 <= U45_in;
    U8 <= U46_in;
    U9 <= U47_in;

    X <= X30_in;

    Y1 <= Y13_in;
    Y2 <= Y14_in;
    Y3 <= Y15_in;
    Y4 <= Y29_in;
    Y5 <= Y30_in;
    Y6 <= Y31_in;
    Y7 <= Y45_in;
    Y8 <= Y46_in;
    Y9 <= Y47_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11110) begin // 31

    Y30_next <= Y_onebyoneout;
    X30_next <= X_onebyoneout;

    U1 <= U14_in;
    U2 <= U15_in;
    U3 <= U16_in;
    U4 <= U30_in;
    U5 <= U31_in;
    U6 <= U32_in;
    U7 <= U46_in;
    U8 <= U47_in;
    U9 <= U48_in;

    X <= X31_in;

    Y1 <= Y14_in;
    Y2 <= Y15_in;
    Y3 <= Y16_in;
    Y4 <= Y30_in;
    Y5 <= Y31_in;
    Y6 <= Y32_in;
    Y7 <= Y46_in;
    Y8 <= Y47_in;
    Y9 <= Y48_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11111) begin // 32

    Y31_next <= Y_onebyoneout;
    X31_next <= X_onebyoneout;

    U1 <= U15_in;
    U2 <= U16_in;
    U3 <= `WIDTH'b0;
    U4 <= U31_in;
    U5 <= U32_in;
    U6 <= `WIDTH'b0;
    U7 <= U47_in;
    U8 <= U48_in;
    U9 <= `WIDTH'b0;

    X <= X32_in;

    Y1 <= Y15_in;
    Y2 <= Y16_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y31_in;
    Y5 <= Y32_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y47_in;
    Y8 <= Y48_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b100000) begin // 33

    Y32_next <= Y_onebyoneout;
    X32_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U17_in;
    U3 <= U18_in;
    U4 <= `WIDTH'b0;
    U5 <= U33_in;
    U6 <= U34_in;
    U7 <= `WIDTH'b0;
    U8 <= U49_in;
    U9 <= U50_in;

    X <= X33_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y17_in;
    Y3 <= Y18_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y33_in;
    Y6 <= Y34_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y49_in;
    Y9 <= Y50_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b100001) begin // 34

    Y33_next <= Y_onebyoneout;
    X33_next <= X_onebyoneout;

    U1 <= U17_in;
    U2 <= U18_in;
    U3 <= U19_in;
    U4 <= U33_in;
    U5 <= U34_in;
    U6 <= U35_in;
    U7 <= U49_in;
    U8 <= U50_in;
    U9 <= U51_in;

    X <= X34_in;

    Y1 <= Y17_in;
    Y2 <= Y18_in;
    Y3 <= Y19_in;
    Y4 <= Y33_in;
    Y5 <= Y34_in;
    Y6 <= Y35_in;
    Y7 <= Y49_in;
    Y8 <= Y50_in;
    Y9 <= Y51_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b100010) begin // 35

    Y34_next <= Y_onebyoneout;
    X34_next <= X_onebyoneout;

    U1 <= U18_in;
    U2 <= U19_in;
    U3 <= U20_in;
    U4 <= U34_in;
    U5 <= U35_in;
    U6 <= U36_in;
    U7 <= U50_in;
    U8 <= U51_in;
    U9 <= U52_in;

    X <= X35_in;

    Y1 <= Y18_in;
    Y2 <= Y19_in;
    Y3 <= Y20_in;
    Y4 <= Y34_in;
    Y5 <= Y35_in;
    Y6 <= Y36_in;
    Y7 <= Y50_in;
    Y8 <= Y51_in;
    Y9 <= Y52_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b100011) begin // 36

    Y35_next <= Y_onebyoneout;
    X35_next <= X_onebyoneout;

    U1 <= U19_in;
    U2 <= U20_in;
    U3 <= U21_in;
    U4 <= U35_in;
    U5 <= U36_in;
    U6 <= U37_in;
    U7 <= U51_in;
    U8 <= U52_in;
    U9 <= U53_in;

    X <= X36_in;

    Y1 <= Y19_in;
    Y2 <= Y20_in;
    Y3 <= Y21_in;
    Y4 <= Y35_in;
    Y5 <= Y36_in;
    Y6 <= Y37_in;
    Y7 <= Y51_in;
    Y8 <= Y52_in;
    Y9 <= Y53_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b100100) begin // 37

    Y36_next <= Y_onebyoneout;
    X36_next <= X_onebyoneout;

    U1 <= U20_in;
    U2 <= U21_in;
    U3 <= U22_in;
    U4 <= U36_in;
    U5 <= U37_in;
    U6 <= U38_in;
    U7 <= U52_in;
    U8 <= U53_in;
    U9 <= U54_in;

    X <= X37_in;

    Y1 <= Y20_in;
    Y2 <= Y21_in;
    Y3 <= Y22_in;
    Y4 <= Y36_in;
    Y5 <= Y37_in;
    Y6 <= Y38_in;
    Y7 <= Y52_in;
    Y8 <= Y53_in;
    Y9 <= Y54_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b100101) begin // 38

    Y37_next <= Y_onebyoneout;
    X37_next <= X_onebyoneout;

    U1 <= U21_in;
    U2 <= U22_in;
    U3 <= U23_in;
    U4 <= U37_in;
    U5 <= U38_in;
    U6 <= U39_in;
    U7 <= U53_in;
    U8 <= U54_in;
    U9 <= U55_in;

    X <= X38_in;

    Y1 <= Y21_in;
    Y2 <= Y22_in;
    Y3 <= Y23_in;
    Y4 <= Y37_in;
    Y5 <= Y38_in;
    Y6 <= Y39_in;
    Y7 <= Y53_in;
    Y8 <= Y54_in;
    Y9 <= Y55_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b100110) begin // 39

    Y38_next <= Y_onebyoneout;
    X38_next <= X_onebyoneout;

    U1 <= U22_in;
    U2 <= U23_in;
    U3 <= U24_in;
    U4 <= U38_in;
    U5 <= U39_in;
    U6 <= U40_in;
    U7 <= U54_in;
    U8 <= U55_in;
    U9 <= U56_in;

    X <= X39_in;

    Y1 <= Y22_in;
    Y2 <= Y23_in;
    Y3 <= Y24_in;
    Y4 <= Y38_in;
    Y5 <= Y39_in;
    Y6 <= Y40_in;
    Y7 <= Y54_in;
    Y8 <= Y55_in;
    Y9 <= Y56_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b100111) begin // 40

    Y39_next <= Y_onebyoneout;
    X39_next <= X_onebyoneout;

    U1 <= U23_in;
    U2 <= U24_in;
    U3 <= U25_in;
    U4 <= U39_in;
    U5 <= U40_in;
    U6 <= U41_in;
    U7 <= U55_in;
    U8 <= U56_in;
    U9 <= U57_in;

    X <= X40_in;

    Y1 <= Y23_in;
    Y2 <= Y24_in;
    Y3 <= Y25_in;
    Y4 <= Y39_in;
    Y5 <= Y40_in;
    Y6 <= Y41_in;
    Y7 <= Y55_in;
    Y8 <= Y56_in;
    Y9 <= Y57_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b101000) begin // 41

    Y40_next <= Y_onebyoneout;
    X40_next <= X_onebyoneout;

    U1 <= U24_in;
    U2 <= U25_in;
    U3 <= U26_in;
    U4 <= U40_in;
    U5 <= U41_in;
    U6 <= U42_in;
    U7 <= U56_in;
    U8 <= U57_in;
    U9 <= U58_in;

    X <= X41_in;

    Y1 <= Y24_in;
    Y2 <= Y25_in;
    Y3 <= Y26_in;
    Y4 <= Y40_in;
    Y5 <= Y41_in;
    Y6 <= Y42_in;
    Y7 <= Y56_in;
    Y8 <= Y57_in;
    Y9 <= Y58_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b101001) begin // 42

    Y41_next <= Y_onebyoneout;
    X41_next <= X_onebyoneout;

    U1 <= U25_in;
    U2 <= U26_in;
    U3 <= U27_in;
    U4 <= U41_in;
    U5 <= U42_in;
    U6 <= U43_in;
    U7 <= U57_in;
    U8 <= U58_in;
    U9 <= U59_in;

    X <= X42_in;

    Y1 <= Y25_in;
    Y2 <= Y26_in;
    Y3 <= Y27_in;
    Y4 <= Y41_in;
    Y5 <= Y42_in;
    Y6 <= Y43_in;
    Y7 <= Y57_in;
    Y8 <= Y58_in;
    Y9 <= Y59_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b101010) begin // 43

    Y42_next <= Y_onebyoneout;
    X42_next <= X_onebyoneout;

    U1 <= U26_in;
    U2 <= U27_in;
    U3 <= U28_in;
    U4 <= U42_in;
    U5 <= U43_in;
    U6 <= U44_in;
    U7 <= U58_in;
    U8 <= U59_in;
    U9 <= U60_in;

    X <= X43_in;

    Y1 <= Y26_in;
    Y2 <= Y27_in;
    Y3 <= Y28_in;
    Y4 <= Y42_in;
    Y5 <= Y43_in;
    Y6 <= Y44_in;
    Y7 <= Y58_in;
    Y8 <= Y59_in;
    Y9 <= Y60_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b101011) begin // 44

    Y43_next <= Y_onebyoneout;
    X43_next <= X_onebyoneout;

    U1 <= U27_in;
    U2 <= U28_in;
    U3 <= U29_in;
    U4 <= U43_in;
    U5 <= U44_in;
    U6 <= U45_in;
    U7 <= U59_in;
    U8 <= U60_in;
    U9 <= U61_in;

    X <= X44_in;

    Y1 <= Y27_in;
    Y2 <= Y28_in;
    Y3 <= Y29_in;
    Y4 <= Y43_in;
    Y5 <= Y44_in;
    Y6 <= Y45_in;
    Y7 <= Y59_in;
    Y8 <= Y60_in;
    Y9 <= Y61_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b101100) begin // 45

    Y44_next <= Y_onebyoneout;
    X44_next <= X_onebyoneout;

    U1 <= U28_in;
    U2 <= U29_in;
    U3 <= U30_in;
    U4 <= U44_in;
    U5 <= U45_in;
    U6 <= U46_in;
    U7 <= U60_in;
    U8 <= U61_in;
    U9 <= U62_in;

    X <= X45_in;

    Y1 <= Y28_in;
    Y2 <= Y29_in;
    Y3 <= Y30_in;
    Y4 <= Y44_in;
    Y5 <= Y45_in;
    Y6 <= Y46_in;
    Y7 <= Y60_in;
    Y8 <= Y61_in;
    Y9 <= Y62_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b101101) begin // 46

    Y45_next <= Y_onebyoneout;
    X45_next <= X_onebyoneout;

    U1 <= U29_in;
    U2 <= U30_in;
    U3 <= U31_in;
    U4 <= U45_in;
    U5 <= U46_in;
    U6 <= U47_in;
    U7 <= U61_in;
    U8 <= U62_in;
    U9 <= U63_in;

    X <= X46_in;

    Y1 <= Y29_in;
    Y2 <= Y30_in;
    Y3 <= Y31_in;
    Y4 <= Y45_in;
    Y5 <= Y46_in;
    Y6 <= Y47_in;
    Y7 <= Y61_in;
    Y8 <= Y62_in;
    Y9 <= Y63_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b101110) begin // 47

    Y46_next <= Y_onebyoneout;
    X46_next <= X_onebyoneout;

    U1 <= U30_in;
    U2 <= U31_in;
    U3 <= U32_in;
    U4 <= U46_in;
    U5 <= U47_in;
    U6 <= U48_in;
    U7 <= U62_in;
    U8 <= U63_in;
    U9 <= U64_in;

    X <= X47_in;

    Y1 <= Y30_in;
    Y2 <= Y31_in;
    Y3 <= Y32_in;
    Y4 <= Y46_in;
    Y5 <= Y47_in;
    Y6 <= Y48_in;
    Y7 <= Y62_in;
    Y8 <= Y63_in;
    Y9 <= Y64_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b101111) begin // 48

    Y47_next <= Y_onebyoneout;
    X47_next <= X_onebyoneout;

    U1 <= U31_in;
    U2 <= U32_in;
    U3 <= `WIDTH'b0;
    U4 <= U47_in;
    U5 <= U48_in;
    U6 <= `WIDTH'b0;
    U7 <= U63_in;
    U8 <= U64_in;
    U9 <= `WIDTH'b0;

    X <= X48_in;

    Y1 <= Y31_in;
    Y2 <= Y32_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y47_in;
    Y5 <= Y48_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y63_in;
    Y8 <= Y64_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b110000) begin // 49

    Y48_next <= Y_onebyoneout;
    X48_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U33_in;
    U3 <= U34_in;
    U4 <= `WIDTH'b0;
    U5 <= U49_in;
    U6 <= U50_in;
    U7 <= `WIDTH'b0;
    U8 <= U65_in;
    U9 <= U66_in;

    X <= X49_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y33_in;
    Y3 <= Y34_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y49_in;
    Y6 <= Y50_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y65_in;
    Y9 <= Y66_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b110001) begin // 50

    Y49_next <= Y_onebyoneout;
    X49_next <= X_onebyoneout;

    U1 <= U33_in;
    U2 <= U34_in;
    U3 <= U35_in;
    U4 <= U49_in;
    U5 <= U50_in;
    U6 <= U51_in;
    U7 <= U65_in;
    U8 <= U66_in;
    U9 <= U67_in;

    X <= X50_in;

    Y1 <= Y33_in;
    Y2 <= Y34_in;
    Y3 <= Y35_in;
    Y4 <= Y49_in;
    Y5 <= Y50_in;
    Y6 <= Y51_in;
    Y7 <= Y65_in;
    Y8 <= Y66_in;
    Y9 <= Y67_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b110010) begin // 51

    Y50_next <= Y_onebyoneout;
    X50_next <= X_onebyoneout;

    U1 <= U34_in;
    U2 <= U35_in;
    U3 <= U36_in;
    U4 <= U50_in;
    U5 <= U51_in;
    U6 <= U52_in;
    U7 <= U66_in;
    U8 <= U67_in;
    U9 <= U68_in;

    X <= X51_in;

    Y1 <= Y34_in;
    Y2 <= Y35_in;
    Y3 <= Y36_in;
    Y4 <= Y50_in;
    Y5 <= Y51_in;
    Y6 <= Y52_in;
    Y7 <= Y66_in;
    Y8 <= Y67_in;
    Y9 <= Y68_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b110011) begin // 52

    Y51_next <= Y_onebyoneout;
    X51_next <= X_onebyoneout;

    U1 <= U35_in;
    U2 <= U36_in;
    U3 <= U37_in;
    U4 <= U51_in;
    U5 <= U52_in;
    U6 <= U53_in;
    U7 <= U67_in;
    U8 <= U68_in;
    U9 <= U69_in;

    X <= X52_in;

    Y1 <= Y35_in;
    Y2 <= Y36_in;
    Y3 <= Y37_in;
    Y4 <= Y51_in;
    Y5 <= Y52_in;
    Y6 <= Y53_in;
    Y7 <= Y67_in;
    Y8 <= Y68_in;
    Y9 <= Y69_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b110100) begin // 53

    Y52_next <= Y_onebyoneout;
    X52_next <= X_onebyoneout;

    U1 <= U36_in;
    U2 <= U37_in;
    U3 <= U38_in;
    U4 <= U52_in;
    U5 <= U53_in;
    U6 <= U54_in;
    U7 <= U68_in;
    U8 <= U69_in;
    U9 <= U70_in;

    X <= X53_in;

    Y1 <= Y36_in;
    Y2 <= Y37_in;
    Y3 <= Y38_in;
    Y4 <= Y52_in;
    Y5 <= Y53_in;
    Y6 <= Y54_in;
    Y7 <= Y68_in;
    Y8 <= Y69_in;
    Y9 <= Y70_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b110101) begin // 54

    Y53_next <= Y_onebyoneout;
    X53_next <= X_onebyoneout;

    U1 <= U37_in;
    U2 <= U38_in;
    U3 <= U39_in;
    U4 <= U53_in;
    U5 <= U54_in;
    U6 <= U55_in;
    U7 <= U69_in;
    U8 <= U70_in;
    U9 <= U71_in;

    X <= X54_in;

    Y1 <= Y37_in;
    Y2 <= Y38_in;
    Y3 <= Y39_in;
    Y4 <= Y53_in;
    Y5 <= Y54_in;
    Y6 <= Y55_in;
    Y7 <= Y69_in;
    Y8 <= Y70_in;
    Y9 <= Y71_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b110110) begin // 55

    Y54_next <= Y_onebyoneout;
    X54_next <= X_onebyoneout;

    U1 <= U38_in;
    U2 <= U39_in;
    U3 <= U40_in;
    U4 <= U54_in;
    U5 <= U55_in;
    U6 <= U56_in;
    U7 <= U70_in;
    U8 <= U71_in;
    U9 <= U72_in;

    X <= X55_in;

    Y1 <= Y38_in;
    Y2 <= Y39_in;
    Y3 <= Y40_in;
    Y4 <= Y54_in;
    Y5 <= Y55_in;
    Y6 <= Y56_in;
    Y7 <= Y70_in;
    Y8 <= Y71_in;
    Y9 <= Y72_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b110111) begin // 56

    Y55_next <= Y_onebyoneout;
    X55_next <= X_onebyoneout;

    U1 <= U39_in;
    U2 <= U40_in;
    U3 <= U41_in;
    U4 <= U55_in;
    U5 <= U56_in;
    U6 <= U57_in;
    U7 <= U71_in;
    U8 <= U72_in;
    U9 <= U73_in;

    X <= X56_in;

    Y1 <= Y39_in;
    Y2 <= Y40_in;
    Y3 <= Y41_in;
    Y4 <= Y55_in;
    Y5 <= Y56_in;
    Y6 <= Y57_in;
    Y7 <= Y71_in;
    Y8 <= Y72_in;
    Y9 <= Y73_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b111000) begin // 57

    Y56_next <= Y_onebyoneout;
    X56_next <= X_onebyoneout;

    U1 <= U40_in;
    U2 <= U41_in;
    U3 <= U42_in;
    U4 <= U56_in;
    U5 <= U57_in;
    U6 <= U58_in;
    U7 <= U72_in;
    U8 <= U73_in;
    U9 <= U74_in;

    X <= X57_in;

    Y1 <= Y40_in;
    Y2 <= Y41_in;
    Y3 <= Y42_in;
    Y4 <= Y56_in;
    Y5 <= Y57_in;
    Y6 <= Y58_in;
    Y7 <= Y72_in;
    Y8 <= Y73_in;
    Y9 <= Y74_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b111001) begin // 58

    Y57_next <= Y_onebyoneout;
    X57_next <= X_onebyoneout;

    U1 <= U41_in;
    U2 <= U42_in;
    U3 <= U43_in;
    U4 <= U57_in;
    U5 <= U58_in;
    U6 <= U59_in;
    U7 <= U73_in;
    U8 <= U74_in;
    U9 <= U75_in;

    X <= X58_in;

    Y1 <= Y41_in;
    Y2 <= Y42_in;
    Y3 <= Y43_in;
    Y4 <= Y57_in;
    Y5 <= Y58_in;
    Y6 <= Y59_in;
    Y7 <= Y73_in;
    Y8 <= Y74_in;
    Y9 <= Y75_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b111010) begin // 59

    Y58_next <= Y_onebyoneout;
    X58_next <= X_onebyoneout;

    U1 <= U42_in;
    U2 <= U43_in;
    U3 <= U44_in;
    U4 <= U58_in;
    U5 <= U59_in;
    U6 <= U60_in;
    U7 <= U74_in;
    U8 <= U75_in;
    U9 <= U76_in;

    X <= X59_in;

    Y1 <= Y42_in;
    Y2 <= Y43_in;
    Y3 <= Y44_in;
    Y4 <= Y58_in;
    Y5 <= Y59_in;
    Y6 <= Y60_in;
    Y7 <= Y74_in;
    Y8 <= Y75_in;
    Y9 <= Y76_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b111011) begin // 60

    Y59_next <= Y_onebyoneout;
    X59_next <= X_onebyoneout;

    U1 <= U43_in;
    U2 <= U44_in;
    U3 <= U45_in;
    U4 <= U59_in;
    U5 <= U60_in;
    U6 <= U61_in;
    U7 <= U75_in;
    U8 <= U76_in;
    U9 <= U77_in;

    X <= X60_in;

    Y1 <= Y43_in;
    Y2 <= Y44_in;
    Y3 <= Y45_in;
    Y4 <= Y59_in;
    Y5 <= Y60_in;
    Y6 <= Y61_in;
    Y7 <= Y75_in;
    Y8 <= Y76_in;
    Y9 <= Y77_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b111100) begin // 61

    Y60_next <= Y_onebyoneout;
    X60_next <= X_onebyoneout;

    U1 <= U44_in;
    U2 <= U45_in;
    U3 <= U46_in;
    U4 <= U60_in;
    U5 <= U61_in;
    U6 <= U62_in;
    U7 <= U76_in;
    U8 <= U77_in;
    U9 <= U78_in;

    X <= X61_in;

    Y1 <= Y44_in;
    Y2 <= Y45_in;
    Y3 <= Y46_in;
    Y4 <= Y60_in;
    Y5 <= Y61_in;
    Y6 <= Y62_in;
    Y7 <= Y76_in;
    Y8 <= Y77_in;
    Y9 <= Y78_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b111101) begin // 62

    Y61_next <= Y_onebyoneout;
    X61_next <= X_onebyoneout;

    U1 <= U45_in;
    U2 <= U46_in;
    U3 <= U47_in;
    U4 <= U61_in;
    U5 <= U62_in;
    U6 <= U63_in;
    U7 <= U77_in;
    U8 <= U78_in;
    U9 <= U79_in;

    X <= X62_in;

    Y1 <= Y45_in;
    Y2 <= Y46_in;
    Y3 <= Y47_in;
    Y4 <= Y61_in;
    Y5 <= Y62_in;
    Y6 <= Y63_in;
    Y7 <= Y77_in;
    Y8 <= Y78_in;
    Y9 <= Y79_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b111110) begin // 63

    Y62_next <= Y_onebyoneout;
    X62_next <= X_onebyoneout;

    U1 <= U46_in;
    U2 <= U47_in;
    U3 <= U48_in;
    U4 <= U62_in;
    U5 <= U63_in;
    U6 <= U64_in;
    U7 <= U78_in;
    U8 <= U79_in;
    U9 <= U80_in;

    X <= X63_in;

    Y1 <= Y46_in;
    Y2 <= Y47_in;
    Y3 <= Y48_in;
    Y4 <= Y62_in;
    Y5 <= Y63_in;
    Y6 <= Y64_in;
    Y7 <= Y78_in;
    Y8 <= Y79_in;
    Y9 <= Y80_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b111111) begin // 64

    Y63_next <= Y_onebyoneout;
    X63_next <= X_onebyoneout;

    U1 <= U47_in;
    U2 <= U48_in;
    U3 <= `WIDTH'b0;
    U4 <= U63_in;
    U5 <= U64_in;
    U6 <= `WIDTH'b0;
    U7 <= U79_in;
    U8 <= U80_in;
    U9 <= `WIDTH'b0;

    X <= X64_in;

    Y1 <= Y47_in;
    Y2 <= Y48_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y63_in;
    Y5 <= Y64_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y79_in;
    Y8 <= Y80_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1000000) begin // 65

    Y64_next <= Y_onebyoneout;
    X64_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U49_in;
    U3 <= U50_in;
    U4 <= `WIDTH'b0;
    U5 <= U65_in;
    U6 <= U66_in;
    U7 <= `WIDTH'b0;
    U8 <= U81_in;
    U9 <= U82_in;

    X <= X65_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y49_in;
    Y3 <= Y50_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y65_in;
    Y6 <= Y66_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y81_in;
    Y9 <= Y82_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1000001) begin // 66

    Y65_next <= Y_onebyoneout;
    X65_next <= X_onebyoneout;

    U1 <= U49_in;
    U2 <= U50_in;
    U3 <= U51_in;
    U4 <= U65_in;
    U5 <= U66_in;
    U6 <= U67_in;
    U7 <= U81_in;
    U8 <= U82_in;
    U9 <= U83_in;

    X <= X66_in;

    Y1 <= Y49_in;
    Y2 <= Y50_in;
    Y3 <= Y51_in;
    Y4 <= Y65_in;
    Y5 <= Y66_in;
    Y6 <= Y67_in;
    Y7 <= Y81_in;
    Y8 <= Y82_in;
    Y9 <= Y83_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1000010) begin // 67

    Y66_next <= Y_onebyoneout;
    X66_next <= X_onebyoneout;

    U1 <= U50_in;
    U2 <= U51_in;
    U3 <= U52_in;
    U4 <= U66_in;
    U5 <= U67_in;
    U6 <= U68_in;
    U7 <= U82_in;
    U8 <= U83_in;
    U9 <= U84_in;

    X <= X67_in;

    Y1 <= Y50_in;
    Y2 <= Y51_in;
    Y3 <= Y52_in;
    Y4 <= Y66_in;
    Y5 <= Y67_in;
    Y6 <= Y68_in;
    Y7 <= Y82_in;
    Y8 <= Y83_in;
    Y9 <= Y84_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1000011) begin // 68

    Y67_next <= Y_onebyoneout;
    X67_next <= X_onebyoneout;

    U1 <= U51_in;
    U2 <= U52_in;
    U3 <= U53_in;
    U4 <= U67_in;
    U5 <= U68_in;
    U6 <= U69_in;
    U7 <= U83_in;
    U8 <= U84_in;
    U9 <= U85_in;

    X <= X68_in;

    Y1 <= Y51_in;
    Y2 <= Y52_in;
    Y3 <= Y53_in;
    Y4 <= Y67_in;
    Y5 <= Y68_in;
    Y6 <= Y69_in;
    Y7 <= Y83_in;
    Y8 <= Y84_in;
    Y9 <= Y85_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1000100) begin // 69

    Y68_next <= Y_onebyoneout;
    X68_next <= X_onebyoneout;

    U1 <= U52_in;
    U2 <= U53_in;
    U3 <= U54_in;
    U4 <= U68_in;
    U5 <= U69_in;
    U6 <= U70_in;
    U7 <= U84_in;
    U8 <= U85_in;
    U9 <= U86_in;

    X <= X69_in;

    Y1 <= Y52_in;
    Y2 <= Y53_in;
    Y3 <= Y54_in;
    Y4 <= Y68_in;
    Y5 <= Y69_in;
    Y6 <= Y70_in;
    Y7 <= Y84_in;
    Y8 <= Y85_in;
    Y9 <= Y86_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1000101) begin // 70

    Y69_next <= Y_onebyoneout;
    X69_next <= X_onebyoneout;

    U1 <= U53_in;
    U2 <= U54_in;
    U3 <= U55_in;
    U4 <= U69_in;
    U5 <= U70_in;
    U6 <= U71_in;
    U7 <= U85_in;
    U8 <= U86_in;
    U9 <= U87_in;

    X <= X70_in;

    Y1 <= Y53_in;
    Y2 <= Y54_in;
    Y3 <= Y55_in;
    Y4 <= Y69_in;
    Y5 <= Y70_in;
    Y6 <= Y71_in;
    Y7 <= Y85_in;
    Y8 <= Y86_in;
    Y9 <= Y87_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1000110) begin // 71

    Y70_next <= Y_onebyoneout;
    X70_next <= X_onebyoneout;

    U1 <= U54_in;
    U2 <= U55_in;
    U3 <= U56_in;
    U4 <= U70_in;
    U5 <= U71_in;
    U6 <= U72_in;
    U7 <= U86_in;
    U8 <= U87_in;
    U9 <= U88_in;

    X <= X71_in;

    Y1 <= Y54_in;
    Y2 <= Y55_in;
    Y3 <= Y56_in;
    Y4 <= Y70_in;
    Y5 <= Y71_in;
    Y6 <= Y72_in;
    Y7 <= Y86_in;
    Y8 <= Y87_in;
    Y9 <= Y88_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1000111) begin // 72

    Y71_next <= Y_onebyoneout;
    X71_next <= X_onebyoneout;

    U1 <= U55_in;
    U2 <= U56_in;
    U3 <= U57_in;
    U4 <= U71_in;
    U5 <= U72_in;
    U6 <= U73_in;
    U7 <= U87_in;
    U8 <= U88_in;
    U9 <= U89_in;

    X <= X72_in;

    Y1 <= Y55_in;
    Y2 <= Y56_in;
    Y3 <= Y57_in;
    Y4 <= Y71_in;
    Y5 <= Y72_in;
    Y6 <= Y73_in;
    Y7 <= Y87_in;
    Y8 <= Y88_in;
    Y9 <= Y89_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1001000) begin // 73

    Y72_next <= Y_onebyoneout;
    X72_next <= X_onebyoneout;

    U1 <= U56_in;
    U2 <= U57_in;
    U3 <= U58_in;
    U4 <= U72_in;
    U5 <= U73_in;
    U6 <= U74_in;
    U7 <= U88_in;
    U8 <= U89_in;
    U9 <= U90_in;

    X <= X73_in;

    Y1 <= Y56_in;
    Y2 <= Y57_in;
    Y3 <= Y58_in;
    Y4 <= Y72_in;
    Y5 <= Y73_in;
    Y6 <= Y74_in;
    Y7 <= Y88_in;
    Y8 <= Y89_in;
    Y9 <= Y90_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1001001) begin // 74

    Y73_next <= Y_onebyoneout;
    X73_next <= X_onebyoneout;

    U1 <= U57_in;
    U2 <= U58_in;
    U3 <= U59_in;
    U4 <= U73_in;
    U5 <= U74_in;
    U6 <= U75_in;
    U7 <= U89_in;
    U8 <= U90_in;
    U9 <= U91_in;

    X <= X74_in;

    Y1 <= Y57_in;
    Y2 <= Y58_in;
    Y3 <= Y59_in;
    Y4 <= Y73_in;
    Y5 <= Y74_in;
    Y6 <= Y75_in;
    Y7 <= Y89_in;
    Y8 <= Y90_in;
    Y9 <= Y91_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1001010) begin // 75

    Y74_next <= Y_onebyoneout;
    X74_next <= X_onebyoneout;

    U1 <= U58_in;
    U2 <= U59_in;
    U3 <= U60_in;
    U4 <= U74_in;
    U5 <= U75_in;
    U6 <= U76_in;
    U7 <= U90_in;
    U8 <= U91_in;
    U9 <= U92_in;

    X <= X75_in;

    Y1 <= Y58_in;
    Y2 <= Y59_in;
    Y3 <= Y60_in;
    Y4 <= Y74_in;
    Y5 <= Y75_in;
    Y6 <= Y76_in;
    Y7 <= Y90_in;
    Y8 <= Y91_in;
    Y9 <= Y92_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1001011) begin // 76

    Y75_next <= Y_onebyoneout;
    X75_next <= X_onebyoneout;

    U1 <= U59_in;
    U2 <= U60_in;
    U3 <= U61_in;
    U4 <= U75_in;
    U5 <= U76_in;
    U6 <= U77_in;
    U7 <= U91_in;
    U8 <= U92_in;
    U9 <= U93_in;

    X <= X76_in;

    Y1 <= Y59_in;
    Y2 <= Y60_in;
    Y3 <= Y61_in;
    Y4 <= Y75_in;
    Y5 <= Y76_in;
    Y6 <= Y77_in;
    Y7 <= Y91_in;
    Y8 <= Y92_in;
    Y9 <= Y93_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1001100) begin // 77

    Y76_next <= Y_onebyoneout;
    X76_next <= X_onebyoneout;

    U1 <= U60_in;
    U2 <= U61_in;
    U3 <= U62_in;
    U4 <= U76_in;
    U5 <= U77_in;
    U6 <= U78_in;
    U7 <= U92_in;
    U8 <= U93_in;
    U9 <= U94_in;

    X <= X77_in;

    Y1 <= Y60_in;
    Y2 <= Y61_in;
    Y3 <= Y62_in;
    Y4 <= Y76_in;
    Y5 <= Y77_in;
    Y6 <= Y78_in;
    Y7 <= Y92_in;
    Y8 <= Y93_in;
    Y9 <= Y94_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1001101) begin // 78

    Y77_next <= Y_onebyoneout;
    X77_next <= X_onebyoneout;

    U1 <= U61_in;
    U2 <= U62_in;
    U3 <= U63_in;
    U4 <= U77_in;
    U5 <= U78_in;
    U6 <= U79_in;
    U7 <= U93_in;
    U8 <= U94_in;
    U9 <= U95_in;

    X <= X78_in;

    Y1 <= Y61_in;
    Y2 <= Y62_in;
    Y3 <= Y63_in;
    Y4 <= Y77_in;
    Y5 <= Y78_in;
    Y6 <= Y79_in;
    Y7 <= Y93_in;
    Y8 <= Y94_in;
    Y9 <= Y95_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1001110) begin // 79

    Y78_next <= Y_onebyoneout;
    X78_next <= X_onebyoneout;

    U1 <= U62_in;
    U2 <= U63_in;
    U3 <= U64_in;
    U4 <= U78_in;
    U5 <= U79_in;
    U6 <= U80_in;
    U7 <= U94_in;
    U8 <= U95_in;
    U9 <= U96_in;

    X <= X79_in;

    Y1 <= Y62_in;
    Y2 <= Y63_in;
    Y3 <= Y64_in;
    Y4 <= Y78_in;
    Y5 <= Y79_in;
    Y6 <= Y80_in;
    Y7 <= Y94_in;
    Y8 <= Y95_in;
    Y9 <= Y96_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1001111) begin // 80

    Y79_next <= Y_onebyoneout;
    X79_next <= X_onebyoneout;

    U1 <= U63_in;
    U2 <= U64_in;
    U3 <= `WIDTH'b0;
    U4 <= U79_in;
    U5 <= U80_in;
    U6 <= `WIDTH'b0;
    U7 <= U95_in;
    U8 <= U96_in;
    U9 <= `WIDTH'b0;

    X <= X80_in;

    Y1 <= Y63_in;
    Y2 <= Y64_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y79_in;
    Y5 <= Y80_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y95_in;
    Y8 <= Y96_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1010000) begin // 81

    Y80_next <= Y_onebyoneout;
    X80_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U65_in;
    U3 <= U66_in;
    U4 <= `WIDTH'b0;
    U5 <= U81_in;
    U6 <= U82_in;
    U7 <= `WIDTH'b0;
    U8 <= U97_in;
    U9 <= U98_in;

    X <= X81_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y65_in;
    Y3 <= Y66_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y81_in;
    Y6 <= Y82_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y97_in;
    Y9 <= Y98_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1010001) begin // 82

    Y81_next <= Y_onebyoneout;
    X81_next <= X_onebyoneout;

    U1 <= U65_in;
    U2 <= U66_in;
    U3 <= U67_in;
    U4 <= U81_in;
    U5 <= U82_in;
    U6 <= U83_in;
    U7 <= U97_in;
    U8 <= U98_in;
    U9 <= U99_in;

    X <= X82_in;

    Y1 <= Y65_in;
    Y2 <= Y66_in;
    Y3 <= Y67_in;
    Y4 <= Y81_in;
    Y5 <= Y82_in;
    Y6 <= Y83_in;
    Y7 <= Y97_in;
    Y8 <= Y98_in;
    Y9 <= Y99_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1010010) begin // 83

    Y82_next <= Y_onebyoneout;
    X82_next <= X_onebyoneout;

    U1 <= U66_in;
    U2 <= U67_in;
    U3 <= U68_in;
    U4 <= U82_in;
    U5 <= U83_in;
    U6 <= U84_in;
    U7 <= U98_in;
    U8 <= U99_in;
    U9 <= U100_in;

    X <= X83_in;

    Y1 <= Y66_in;
    Y2 <= Y67_in;
    Y3 <= Y68_in;
    Y4 <= Y82_in;
    Y5 <= Y83_in;
    Y6 <= Y84_in;
    Y7 <= Y98_in;
    Y8 <= Y99_in;
    Y9 <= Y100_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1010011) begin // 84

    Y83_next <= Y_onebyoneout;
    X83_next <= X_onebyoneout;

    U1 <= U67_in;
    U2 <= U68_in;
    U3 <= U69_in;
    U4 <= U83_in;
    U5 <= U84_in;
    U6 <= U85_in;
    U7 <= U99_in;
    U8 <= U100_in;
    U9 <= U101_in;

    X <= X84_in;

    Y1 <= Y67_in;
    Y2 <= Y68_in;
    Y3 <= Y69_in;
    Y4 <= Y83_in;
    Y5 <= Y84_in;
    Y6 <= Y85_in;
    Y7 <= Y99_in;
    Y8 <= Y100_in;
    Y9 <= Y101_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1010100) begin // 85

    Y84_next <= Y_onebyoneout;
    X84_next <= X_onebyoneout;

    U1 <= U68_in;
    U2 <= U69_in;
    U3 <= U70_in;
    U4 <= U84_in;
    U5 <= U85_in;
    U6 <= U86_in;
    U7 <= U100_in;
    U8 <= U101_in;
    U9 <= U102_in;

    X <= X85_in;

    Y1 <= Y68_in;
    Y2 <= Y69_in;
    Y3 <= Y70_in;
    Y4 <= Y84_in;
    Y5 <= Y85_in;
    Y6 <= Y86_in;
    Y7 <= Y100_in;
    Y8 <= Y101_in;
    Y9 <= Y102_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1010101) begin // 86

    Y85_next <= Y_onebyoneout;
    X85_next <= X_onebyoneout;

    U1 <= U69_in;
    U2 <= U70_in;
    U3 <= U71_in;
    U4 <= U85_in;
    U5 <= U86_in;
    U6 <= U87_in;
    U7 <= U101_in;
    U8 <= U102_in;
    U9 <= U103_in;

    X <= X86_in;

    Y1 <= Y69_in;
    Y2 <= Y70_in;
    Y3 <= Y71_in;
    Y4 <= Y85_in;
    Y5 <= Y86_in;
    Y6 <= Y87_in;
    Y7 <= Y101_in;
    Y8 <= Y102_in;
    Y9 <= Y103_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1010110) begin // 87

    Y86_next <= Y_onebyoneout;
    X86_next <= X_onebyoneout;

    U1 <= U70_in;
    U2 <= U71_in;
    U3 <= U72_in;
    U4 <= U86_in;
    U5 <= U87_in;
    U6 <= U88_in;
    U7 <= U102_in;
    U8 <= U103_in;
    U9 <= U104_in;

    X <= X87_in;

    Y1 <= Y70_in;
    Y2 <= Y71_in;
    Y3 <= Y72_in;
    Y4 <= Y86_in;
    Y5 <= Y87_in;
    Y6 <= Y88_in;
    Y7 <= Y102_in;
    Y8 <= Y103_in;
    Y9 <= Y104_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1010111) begin // 88

    Y87_next <= Y_onebyoneout;
    X87_next <= X_onebyoneout;

    U1 <= U71_in;
    U2 <= U72_in;
    U3 <= U73_in;
    U4 <= U87_in;
    U5 <= U88_in;
    U6 <= U89_in;
    U7 <= U103_in;
    U8 <= U104_in;
    U9 <= U105_in;

    X <= X88_in;

    Y1 <= Y71_in;
    Y2 <= Y72_in;
    Y3 <= Y73_in;
    Y4 <= Y87_in;
    Y5 <= Y88_in;
    Y6 <= Y89_in;
    Y7 <= Y103_in;
    Y8 <= Y104_in;
    Y9 <= Y105_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1011000) begin // 89

    Y88_next <= Y_onebyoneout;
    X88_next <= X_onebyoneout;

    U1 <= U72_in;
    U2 <= U73_in;
    U3 <= U74_in;
    U4 <= U88_in;
    U5 <= U89_in;
    U6 <= U90_in;
    U7 <= U104_in;
    U8 <= U105_in;
    U9 <= U106_in;

    X <= X89_in;

    Y1 <= Y72_in;
    Y2 <= Y73_in;
    Y3 <= Y74_in;
    Y4 <= Y88_in;
    Y5 <= Y89_in;
    Y6 <= Y90_in;
    Y7 <= Y104_in;
    Y8 <= Y105_in;
    Y9 <= Y106_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1011001) begin // 90

    Y89_next <= Y_onebyoneout;
    X89_next <= X_onebyoneout;

    U1 <= U73_in;
    U2 <= U74_in;
    U3 <= U75_in;
    U4 <= U89_in;
    U5 <= U90_in;
    U6 <= U91_in;
    U7 <= U105_in;
    U8 <= U106_in;
    U9 <= U107_in;

    X <= X90_in;

    Y1 <= Y73_in;
    Y2 <= Y74_in;
    Y3 <= Y75_in;
    Y4 <= Y89_in;
    Y5 <= Y90_in;
    Y6 <= Y91_in;
    Y7 <= Y105_in;
    Y8 <= Y106_in;
    Y9 <= Y107_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1011010) begin // 91

    Y90_next <= Y_onebyoneout;
    X90_next <= X_onebyoneout;

    U1 <= U74_in;
    U2 <= U75_in;
    U3 <= U76_in;
    U4 <= U90_in;
    U5 <= U91_in;
    U6 <= U92_in;
    U7 <= U106_in;
    U8 <= U107_in;
    U9 <= U108_in;

    X <= X91_in;

    Y1 <= Y74_in;
    Y2 <= Y75_in;
    Y3 <= Y76_in;
    Y4 <= Y90_in;
    Y5 <= Y91_in;
    Y6 <= Y92_in;
    Y7 <= Y106_in;
    Y8 <= Y107_in;
    Y9 <= Y108_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1011011) begin // 92

    Y91_next <= Y_onebyoneout;
    X91_next <= X_onebyoneout;

    U1 <= U75_in;
    U2 <= U76_in;
    U3 <= U77_in;
    U4 <= U91_in;
    U5 <= U92_in;
    U6 <= U93_in;
    U7 <= U107_in;
    U8 <= U108_in;
    U9 <= U109_in;

    X <= X92_in;

    Y1 <= Y75_in;
    Y2 <= Y76_in;
    Y3 <= Y77_in;
    Y4 <= Y91_in;
    Y5 <= Y92_in;
    Y6 <= Y93_in;
    Y7 <= Y107_in;
    Y8 <= Y108_in;
    Y9 <= Y109_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1011100) begin // 93

    Y92_next <= Y_onebyoneout;
    X92_next <= X_onebyoneout;

    U1 <= U76_in;
    U2 <= U77_in;
    U3 <= U78_in;
    U4 <= U92_in;
    U5 <= U93_in;
    U6 <= U94_in;
    U7 <= U108_in;
    U8 <= U109_in;
    U9 <= U110_in;

    X <= X93_in;

    Y1 <= Y76_in;
    Y2 <= Y77_in;
    Y3 <= Y78_in;
    Y4 <= Y92_in;
    Y5 <= Y93_in;
    Y6 <= Y94_in;
    Y7 <= Y108_in;
    Y8 <= Y109_in;
    Y9 <= Y110_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1011101) begin // 94

    Y93_next <= Y_onebyoneout;
    X93_next <= X_onebyoneout;

    U1 <= U77_in;
    U2 <= U78_in;
    U3 <= U79_in;
    U4 <= U93_in;
    U5 <= U94_in;
    U6 <= U95_in;
    U7 <= U109_in;
    U8 <= U110_in;
    U9 <= U111_in;

    X <= X94_in;

    Y1 <= Y77_in;
    Y2 <= Y78_in;
    Y3 <= Y79_in;
    Y4 <= Y93_in;
    Y5 <= Y94_in;
    Y6 <= Y95_in;
    Y7 <= Y109_in;
    Y8 <= Y110_in;
    Y9 <= Y111_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1011110) begin // 95

    Y94_next <= Y_onebyoneout;
    X94_next <= X_onebyoneout;

    U1 <= U78_in;
    U2 <= U79_in;
    U3 <= U80_in;
    U4 <= U94_in;
    U5 <= U95_in;
    U6 <= U96_in;
    U7 <= U110_in;
    U8 <= U111_in;
    U9 <= U112_in;

    X <= X95_in;

    Y1 <= Y78_in;
    Y2 <= Y79_in;
    Y3 <= Y80_in;
    Y4 <= Y94_in;
    Y5 <= Y95_in;
    Y6 <= Y96_in;
    Y7 <= Y110_in;
    Y8 <= Y111_in;
    Y9 <= Y112_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1011111) begin // 96

    Y95_next <= Y_onebyoneout;
    X95_next <= X_onebyoneout;

    U1 <= U79_in;
    U2 <= U80_in;
    U3 <= `WIDTH'b0;
    U4 <= U95_in;
    U5 <= U96_in;
    U6 <= `WIDTH'b0;
    U7 <= U111_in;
    U8 <= U112_in;
    U9 <= `WIDTH'b0;

    X <= X96_in;

    Y1 <= Y79_in;
    Y2 <= Y80_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y95_in;
    Y5 <= Y96_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y111_in;
    Y8 <= Y112_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1100000) begin // 97

    Y96_next <= Y_onebyoneout;
    X96_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U81_in;
    U3 <= U82_in;
    U4 <= `WIDTH'b0;
    U5 <= U97_in;
    U6 <= U98_in;
    U7 <= `WIDTH'b0;
    U8 <= U113_in;
    U9 <= U114_in;

    X <= X97_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y81_in;
    Y3 <= Y82_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y97_in;
    Y6 <= Y98_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y113_in;
    Y9 <= Y114_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1100001) begin // 98

    Y97_next <= Y_onebyoneout;
    X97_next <= X_onebyoneout;

    U1 <= U81_in;
    U2 <= U82_in;
    U3 <= U83_in;
    U4 <= U97_in;
    U5 <= U98_in;
    U6 <= U99_in;
    U7 <= U113_in;
    U8 <= U114_in;
    U9 <= U115_in;

    X <= X98_in;

    Y1 <= Y81_in;
    Y2 <= Y82_in;
    Y3 <= Y83_in;
    Y4 <= Y97_in;
    Y5 <= Y98_in;
    Y6 <= Y99_in;
    Y7 <= Y113_in;
    Y8 <= Y114_in;
    Y9 <= Y115_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1100010) begin // 99

    Y98_next <= Y_onebyoneout;
    X98_next <= X_onebyoneout;

    U1 <= U82_in;
    U2 <= U83_in;
    U3 <= U84_in;
    U4 <= U98_in;
    U5 <= U99_in;
    U6 <= U100_in;
    U7 <= U114_in;
    U8 <= U115_in;
    U9 <= U116_in;

    X <= X99_in;

    Y1 <= Y82_in;
    Y2 <= Y83_in;
    Y3 <= Y84_in;
    Y4 <= Y98_in;
    Y5 <= Y99_in;
    Y6 <= Y100_in;
    Y7 <= Y114_in;
    Y8 <= Y115_in;
    Y9 <= Y116_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1100011) begin // 100

    Y99_next <= Y_onebyoneout;
    X99_next <= X_onebyoneout;

    U1 <= U83_in;
    U2 <= U84_in;
    U3 <= U85_in;
    U4 <= U99_in;
    U5 <= U100_in;
    U6 <= U101_in;
    U7 <= U115_in;
    U8 <= U116_in;
    U9 <= U117_in;

    X <= X100_in;

    Y1 <= Y83_in;
    Y2 <= Y84_in;
    Y3 <= Y85_in;
    Y4 <= Y99_in;
    Y5 <= Y100_in;
    Y6 <= Y101_in;
    Y7 <= Y115_in;
    Y8 <= Y116_in;
    Y9 <= Y117_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1100100) begin // 101

    Y100_next <= Y_onebyoneout;
    X100_next <= X_onebyoneout;

    U1 <= U84_in;
    U2 <= U85_in;
    U3 <= U86_in;
    U4 <= U100_in;
    U5 <= U101_in;
    U6 <= U102_in;
    U7 <= U116_in;
    U8 <= U117_in;
    U9 <= U118_in;

    X <= X101_in;

    Y1 <= Y84_in;
    Y2 <= Y85_in;
    Y3 <= Y86_in;
    Y4 <= Y100_in;
    Y5 <= Y101_in;
    Y6 <= Y102_in;
    Y7 <= Y116_in;
    Y8 <= Y117_in;
    Y9 <= Y118_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1100101) begin // 102

    Y101_next <= Y_onebyoneout;
    X101_next <= X_onebyoneout;

    U1 <= U85_in;
    U2 <= U86_in;
    U3 <= U87_in;
    U4 <= U101_in;
    U5 <= U102_in;
    U6 <= U103_in;
    U7 <= U117_in;
    U8 <= U118_in;
    U9 <= U119_in;

    X <= X102_in;

    Y1 <= Y85_in;
    Y2 <= Y86_in;
    Y3 <= Y87_in;
    Y4 <= Y101_in;
    Y5 <= Y102_in;
    Y6 <= Y103_in;
    Y7 <= Y117_in;
    Y8 <= Y118_in;
    Y9 <= Y119_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1100110) begin // 103

    Y102_next <= Y_onebyoneout;
    X102_next <= X_onebyoneout;

    U1 <= U86_in;
    U2 <= U87_in;
    U3 <= U88_in;
    U4 <= U102_in;
    U5 <= U103_in;
    U6 <= U104_in;
    U7 <= U118_in;
    U8 <= U119_in;
    U9 <= U120_in;

    X <= X103_in;

    Y1 <= Y86_in;
    Y2 <= Y87_in;
    Y3 <= Y88_in;
    Y4 <= Y102_in;
    Y5 <= Y103_in;
    Y6 <= Y104_in;
    Y7 <= Y118_in;
    Y8 <= Y119_in;
    Y9 <= Y120_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1100111) begin // 104

    Y103_next <= Y_onebyoneout;
    X103_next <= X_onebyoneout;

    U1 <= U87_in;
    U2 <= U88_in;
    U3 <= U89_in;
    U4 <= U103_in;
    U5 <= U104_in;
    U6 <= U105_in;
    U7 <= U119_in;
    U8 <= U120_in;
    U9 <= U121_in;

    X <= X104_in;

    Y1 <= Y87_in;
    Y2 <= Y88_in;
    Y3 <= Y89_in;
    Y4 <= Y103_in;
    Y5 <= Y104_in;
    Y6 <= Y105_in;
    Y7 <= Y119_in;
    Y8 <= Y120_in;
    Y9 <= Y121_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1101000) begin // 105

    Y104_next <= Y_onebyoneout;
    X104_next <= X_onebyoneout;

    U1 <= U88_in;
    U2 <= U89_in;
    U3 <= U90_in;
    U4 <= U104_in;
    U5 <= U105_in;
    U6 <= U106_in;
    U7 <= U120_in;
    U8 <= U121_in;
    U9 <= U122_in;

    X <= X105_in;

    Y1 <= Y88_in;
    Y2 <= Y89_in;
    Y3 <= Y90_in;
    Y4 <= Y104_in;
    Y5 <= Y105_in;
    Y6 <= Y106_in;
    Y7 <= Y120_in;
    Y8 <= Y121_in;
    Y9 <= Y122_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1101001) begin // 106

    Y105_next <= Y_onebyoneout;
    X105_next <= X_onebyoneout;

    U1 <= U89_in;
    U2 <= U90_in;
    U3 <= U91_in;
    U4 <= U105_in;
    U5 <= U106_in;
    U6 <= U107_in;
    U7 <= U121_in;
    U8 <= U122_in;
    U9 <= U123_in;

    X <= X106_in;

    Y1 <= Y89_in;
    Y2 <= Y90_in;
    Y3 <= Y91_in;
    Y4 <= Y105_in;
    Y5 <= Y106_in;
    Y6 <= Y107_in;
    Y7 <= Y121_in;
    Y8 <= Y122_in;
    Y9 <= Y123_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1101010) begin // 107

    Y106_next <= Y_onebyoneout;
    X106_next <= X_onebyoneout;

    U1 <= U90_in;
    U2 <= U91_in;
    U3 <= U92_in;
    U4 <= U106_in;
    U5 <= U107_in;
    U6 <= U108_in;
    U7 <= U122_in;
    U8 <= U123_in;
    U9 <= U124_in;

    X <= X107_in;

    Y1 <= Y90_in;
    Y2 <= Y91_in;
    Y3 <= Y92_in;
    Y4 <= Y106_in;
    Y5 <= Y107_in;
    Y6 <= Y108_in;
    Y7 <= Y122_in;
    Y8 <= Y123_in;
    Y9 <= Y124_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1101011) begin // 108

    Y107_next <= Y_onebyoneout;
    X107_next <= X_onebyoneout;

    U1 <= U91_in;
    U2 <= U92_in;
    U3 <= U93_in;
    U4 <= U107_in;
    U5 <= U108_in;
    U6 <= U109_in;
    U7 <= U123_in;
    U8 <= U124_in;
    U9 <= U125_in;

    X <= X108_in;

    Y1 <= Y91_in;
    Y2 <= Y92_in;
    Y3 <= Y93_in;
    Y4 <= Y107_in;
    Y5 <= Y108_in;
    Y6 <= Y109_in;
    Y7 <= Y123_in;
    Y8 <= Y124_in;
    Y9 <= Y125_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1101100) begin // 109

    Y108_next <= Y_onebyoneout;
    X108_next <= X_onebyoneout;

    U1 <= U92_in;
    U2 <= U93_in;
    U3 <= U94_in;
    U4 <= U108_in;
    U5 <= U109_in;
    U6 <= U110_in;
    U7 <= U124_in;
    U8 <= U125_in;
    U9 <= U126_in;

    X <= X109_in;

    Y1 <= Y92_in;
    Y2 <= Y93_in;
    Y3 <= Y94_in;
    Y4 <= Y108_in;
    Y5 <= Y109_in;
    Y6 <= Y110_in;
    Y7 <= Y124_in;
    Y8 <= Y125_in;
    Y9 <= Y126_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1101101) begin // 110

    Y109_next <= Y_onebyoneout;
    X109_next <= X_onebyoneout;

    U1 <= U93_in;
    U2 <= U94_in;
    U3 <= U95_in;
    U4 <= U109_in;
    U5 <= U110_in;
    U6 <= U111_in;
    U7 <= U125_in;
    U8 <= U126_in;
    U9 <= U127_in;

    X <= X110_in;

    Y1 <= Y93_in;
    Y2 <= Y94_in;
    Y3 <= Y95_in;
    Y4 <= Y109_in;
    Y5 <= Y110_in;
    Y6 <= Y111_in;
    Y7 <= Y125_in;
    Y8 <= Y126_in;
    Y9 <= Y127_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1101110) begin // 111

    Y110_next <= Y_onebyoneout;
    X110_next <= X_onebyoneout;

    U1 <= U94_in;
    U2 <= U95_in;
    U3 <= U96_in;
    U4 <= U110_in;
    U5 <= U111_in;
    U6 <= U112_in;
    U7 <= U126_in;
    U8 <= U127_in;
    U9 <= U128_in;

    X <= X111_in;

    Y1 <= Y94_in;
    Y2 <= Y95_in;
    Y3 <= Y96_in;
    Y4 <= Y110_in;
    Y5 <= Y111_in;
    Y6 <= Y112_in;
    Y7 <= Y126_in;
    Y8 <= Y127_in;
    Y9 <= Y128_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1101111) begin // 112

    Y111_next <= Y_onebyoneout;
    X111_next <= X_onebyoneout;

    U1 <= U95_in;
    U2 <= U96_in;
    U3 <= `WIDTH'b0;
    U4 <= U111_in;
    U5 <= U112_in;
    U6 <= `WIDTH'b0;
    U7 <= U127_in;
    U8 <= U128_in;
    U9 <= `WIDTH'b0;

    X <= X112_in;

    Y1 <= Y95_in;
    Y2 <= Y96_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y111_in;
    Y5 <= Y112_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y127_in;
    Y8 <= Y128_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1110000) begin // 113

    Y112_next <= Y_onebyoneout;
    X112_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U97_in;
    U3 <= U98_in;
    U4 <= `WIDTH'b0;
    U5 <= U113_in;
    U6 <= U114_in;
    U7 <= `WIDTH'b0;
    U8 <= U129_in;
    U9 <= U130_in;

    X <= X113_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y97_in;
    Y3 <= Y98_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y113_in;
    Y6 <= Y114_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y129_in;
    Y9 <= Y130_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1110001) begin // 114

    Y113_next <= Y_onebyoneout;
    X113_next <= X_onebyoneout;

    U1 <= U97_in;
    U2 <= U98_in;
    U3 <= U99_in;
    U4 <= U113_in;
    U5 <= U114_in;
    U6 <= U115_in;
    U7 <= U129_in;
    U8 <= U130_in;
    U9 <= U131_in;

    X <= X114_in;

    Y1 <= Y97_in;
    Y2 <= Y98_in;
    Y3 <= Y99_in;
    Y4 <= Y113_in;
    Y5 <= Y114_in;
    Y6 <= Y115_in;
    Y7 <= Y129_in;
    Y8 <= Y130_in;
    Y9 <= Y131_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1110010) begin // 115

    Y114_next <= Y_onebyoneout;
    X114_next <= X_onebyoneout;

    U1 <= U98_in;
    U2 <= U99_in;
    U3 <= U100_in;
    U4 <= U114_in;
    U5 <= U115_in;
    U6 <= U116_in;
    U7 <= U130_in;
    U8 <= U131_in;
    U9 <= U132_in;

    X <= X115_in;

    Y1 <= Y98_in;
    Y2 <= Y99_in;
    Y3 <= Y100_in;
    Y4 <= Y114_in;
    Y5 <= Y115_in;
    Y6 <= Y116_in;
    Y7 <= Y130_in;
    Y8 <= Y131_in;
    Y9 <= Y132_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1110011) begin // 116

    Y115_next <= Y_onebyoneout;
    X115_next <= X_onebyoneout;

    U1 <= U99_in;
    U2 <= U100_in;
    U3 <= U101_in;
    U4 <= U115_in;
    U5 <= U116_in;
    U6 <= U117_in;
    U7 <= U131_in;
    U8 <= U132_in;
    U9 <= U133_in;

    X <= X116_in;

    Y1 <= Y99_in;
    Y2 <= Y100_in;
    Y3 <= Y101_in;
    Y4 <= Y115_in;
    Y5 <= Y116_in;
    Y6 <= Y117_in;
    Y7 <= Y131_in;
    Y8 <= Y132_in;
    Y9 <= Y133_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1110100) begin // 117

    Y116_next <= Y_onebyoneout;
    X116_next <= X_onebyoneout;

    U1 <= U100_in;
    U2 <= U101_in;
    U3 <= U102_in;
    U4 <= U116_in;
    U5 <= U117_in;
    U6 <= U118_in;
    U7 <= U132_in;
    U8 <= U133_in;
    U9 <= U134_in;

    X <= X117_in;

    Y1 <= Y100_in;
    Y2 <= Y101_in;
    Y3 <= Y102_in;
    Y4 <= Y116_in;
    Y5 <= Y117_in;
    Y6 <= Y118_in;
    Y7 <= Y132_in;
    Y8 <= Y133_in;
    Y9 <= Y134_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1110101) begin // 118

    Y117_next <= Y_onebyoneout;
    X117_next <= X_onebyoneout;

    U1 <= U101_in;
    U2 <= U102_in;
    U3 <= U103_in;
    U4 <= U117_in;
    U5 <= U118_in;
    U6 <= U119_in;
    U7 <= U133_in;
    U8 <= U134_in;
    U9 <= U135_in;

    X <= X118_in;

    Y1 <= Y101_in;
    Y2 <= Y102_in;
    Y3 <= Y103_in;
    Y4 <= Y117_in;
    Y5 <= Y118_in;
    Y6 <= Y119_in;
    Y7 <= Y133_in;
    Y8 <= Y134_in;
    Y9 <= Y135_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1110110) begin // 119

    Y118_next <= Y_onebyoneout;
    X118_next <= X_onebyoneout;

    U1 <= U102_in;
    U2 <= U103_in;
    U3 <= U104_in;
    U4 <= U118_in;
    U5 <= U119_in;
    U6 <= U120_in;
    U7 <= U134_in;
    U8 <= U135_in;
    U9 <= U136_in;

    X <= X119_in;

    Y1 <= Y102_in;
    Y2 <= Y103_in;
    Y3 <= Y104_in;
    Y4 <= Y118_in;
    Y5 <= Y119_in;
    Y6 <= Y120_in;
    Y7 <= Y134_in;
    Y8 <= Y135_in;
    Y9 <= Y136_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1110111) begin // 120

    Y119_next <= Y_onebyoneout;
    X119_next <= X_onebyoneout;

    U1 <= U103_in;
    U2 <= U104_in;
    U3 <= U105_in;
    U4 <= U119_in;
    U5 <= U120_in;
    U6 <= U121_in;
    U7 <= U135_in;
    U8 <= U136_in;
    U9 <= U137_in;

    X <= X120_in;

    Y1 <= Y103_in;
    Y2 <= Y104_in;
    Y3 <= Y105_in;
    Y4 <= Y119_in;
    Y5 <= Y120_in;
    Y6 <= Y121_in;
    Y7 <= Y135_in;
    Y8 <= Y136_in;
    Y9 <= Y137_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1111000) begin // 121

    Y120_next <= Y_onebyoneout;
    X120_next <= X_onebyoneout;

    U1 <= U104_in;
    U2 <= U105_in;
    U3 <= U106_in;
    U4 <= U120_in;
    U5 <= U121_in;
    U6 <= U122_in;
    U7 <= U136_in;
    U8 <= U137_in;
    U9 <= U138_in;

    X <= X121_in;

    Y1 <= Y104_in;
    Y2 <= Y105_in;
    Y3 <= Y106_in;
    Y4 <= Y120_in;
    Y5 <= Y121_in;
    Y6 <= Y122_in;
    Y7 <= Y136_in;
    Y8 <= Y137_in;
    Y9 <= Y138_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1111001) begin // 122

    Y121_next <= Y_onebyoneout;
    X121_next <= X_onebyoneout;

    U1 <= U105_in;
    U2 <= U106_in;
    U3 <= U107_in;
    U4 <= U121_in;
    U5 <= U122_in;
    U6 <= U123_in;
    U7 <= U137_in;
    U8 <= U138_in;
    U9 <= U139_in;

    X <= X122_in;

    Y1 <= Y105_in;
    Y2 <= Y106_in;
    Y3 <= Y107_in;
    Y4 <= Y121_in;
    Y5 <= Y122_in;
    Y6 <= Y123_in;
    Y7 <= Y137_in;
    Y8 <= Y138_in;
    Y9 <= Y139_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1111010) begin // 123

    Y122_next <= Y_onebyoneout;
    X122_next <= X_onebyoneout;

    U1 <= U106_in;
    U2 <= U107_in;
    U3 <= U108_in;
    U4 <= U122_in;
    U5 <= U123_in;
    U6 <= U124_in;
    U7 <= U138_in;
    U8 <= U139_in;
    U9 <= U140_in;

    X <= X123_in;

    Y1 <= Y106_in;
    Y2 <= Y107_in;
    Y3 <= Y108_in;
    Y4 <= Y122_in;
    Y5 <= Y123_in;
    Y6 <= Y124_in;
    Y7 <= Y138_in;
    Y8 <= Y139_in;
    Y9 <= Y140_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1111011) begin // 124

    Y123_next <= Y_onebyoneout;
    X123_next <= X_onebyoneout;

    U1 <= U107_in;
    U2 <= U108_in;
    U3 <= U109_in;
    U4 <= U123_in;
    U5 <= U124_in;
    U6 <= U125_in;
    U7 <= U139_in;
    U8 <= U140_in;
    U9 <= U141_in;

    X <= X124_in;

    Y1 <= Y107_in;
    Y2 <= Y108_in;
    Y3 <= Y109_in;
    Y4 <= Y123_in;
    Y5 <= Y124_in;
    Y6 <= Y125_in;
    Y7 <= Y139_in;
    Y8 <= Y140_in;
    Y9 <= Y141_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1111100) begin // 125

    Y124_next <= Y_onebyoneout;
    X124_next <= X_onebyoneout;

    U1 <= U108_in;
    U2 <= U109_in;
    U3 <= U110_in;
    U4 <= U124_in;
    U5 <= U125_in;
    U6 <= U126_in;
    U7 <= U140_in;
    U8 <= U141_in;
    U9 <= U142_in;

    X <= X125_in;

    Y1 <= Y108_in;
    Y2 <= Y109_in;
    Y3 <= Y110_in;
    Y4 <= Y124_in;
    Y5 <= Y125_in;
    Y6 <= Y126_in;
    Y7 <= Y140_in;
    Y8 <= Y141_in;
    Y9 <= Y142_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1111101) begin // 126

    Y125_next <= Y_onebyoneout;
    X125_next <= X_onebyoneout;

    U1 <= U109_in;
    U2 <= U110_in;
    U3 <= U111_in;
    U4 <= U125_in;
    U5 <= U126_in;
    U6 <= U127_in;
    U7 <= U141_in;
    U8 <= U142_in;
    U9 <= U143_in;

    X <= X126_in;

    Y1 <= Y109_in;
    Y2 <= Y110_in;
    Y3 <= Y111_in;
    Y4 <= Y125_in;
    Y5 <= Y126_in;
    Y6 <= Y127_in;
    Y7 <= Y141_in;
    Y8 <= Y142_in;
    Y9 <= Y143_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1111110) begin // 127

    Y126_next <= Y_onebyoneout;
    X126_next <= X_onebyoneout;

    U1 <= U110_in;
    U2 <= U111_in;
    U3 <= U112_in;
    U4 <= U126_in;
    U5 <= U127_in;
    U6 <= U128_in;
    U7 <= U142_in;
    U8 <= U143_in;
    U9 <= U144_in;

    X <= X127_in;

    Y1 <= Y110_in;
    Y2 <= Y111_in;
    Y3 <= Y112_in;
    Y4 <= Y126_in;
    Y5 <= Y127_in;
    Y6 <= Y128_in;
    Y7 <= Y142_in;
    Y8 <= Y143_in;
    Y9 <= Y144_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1111111) begin // 128

    Y127_next <= Y_onebyoneout;
    X127_next <= X_onebyoneout;

    U1 <= U111_in;
    U2 <= U112_in;
    U3 <= `WIDTH'b0;
    U4 <= U127_in;
    U5 <= U128_in;
    U6 <= `WIDTH'b0;
    U7 <= U143_in;
    U8 <= U144_in;
    U9 <= `WIDTH'b0;

    X <= X128_in;

    Y1 <= Y111_in;
    Y2 <= Y112_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y127_in;
    Y5 <= Y128_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y143_in;
    Y8 <= Y144_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10000000) begin // 129

    Y128_next <= Y_onebyoneout;
    X128_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U113_in;
    U3 <= U114_in;
    U4 <= `WIDTH'b0;
    U5 <= U129_in;
    U6 <= U130_in;
    U7 <= `WIDTH'b0;
    U8 <= U145_in;
    U9 <= U146_in;

    X <= X129_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y113_in;
    Y3 <= Y114_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y129_in;
    Y6 <= Y130_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y145_in;
    Y9 <= Y146_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10000001) begin // 130

    Y129_next <= Y_onebyoneout;
    X129_next <= X_onebyoneout;

    U1 <= U113_in;
    U2 <= U114_in;
    U3 <= U115_in;
    U4 <= U129_in;
    U5 <= U130_in;
    U6 <= U131_in;
    U7 <= U145_in;
    U8 <= U146_in;
    U9 <= U147_in;

    X <= X130_in;

    Y1 <= Y113_in;
    Y2 <= Y114_in;
    Y3 <= Y115_in;
    Y4 <= Y129_in;
    Y5 <= Y130_in;
    Y6 <= Y131_in;
    Y7 <= Y145_in;
    Y8 <= Y146_in;
    Y9 <= Y147_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10000010) begin // 131

    Y130_next <= Y_onebyoneout;
    X130_next <= X_onebyoneout;

    U1 <= U114_in;
    U2 <= U115_in;
    U3 <= U116_in;
    U4 <= U130_in;
    U5 <= U131_in;
    U6 <= U132_in;
    U7 <= U146_in;
    U8 <= U147_in;
    U9 <= U148_in;

    X <= X131_in;

    Y1 <= Y114_in;
    Y2 <= Y115_in;
    Y3 <= Y116_in;
    Y4 <= Y130_in;
    Y5 <= Y131_in;
    Y6 <= Y132_in;
    Y7 <= Y146_in;
    Y8 <= Y147_in;
    Y9 <= Y148_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10000011) begin // 132

    Y131_next <= Y_onebyoneout;
    X131_next <= X_onebyoneout;

    U1 <= U115_in;
    U2 <= U116_in;
    U3 <= U117_in;
    U4 <= U131_in;
    U5 <= U132_in;
    U6 <= U133_in;
    U7 <= U147_in;
    U8 <= U148_in;
    U9 <= U149_in;

    X <= X132_in;

    Y1 <= Y115_in;
    Y2 <= Y116_in;
    Y3 <= Y117_in;
    Y4 <= Y131_in;
    Y5 <= Y132_in;
    Y6 <= Y133_in;
    Y7 <= Y147_in;
    Y8 <= Y148_in;
    Y9 <= Y149_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10000100) begin // 133

    Y132_next <= Y_onebyoneout;
    X132_next <= X_onebyoneout;

    U1 <= U116_in;
    U2 <= U117_in;
    U3 <= U118_in;
    U4 <= U132_in;
    U5 <= U133_in;
    U6 <= U134_in;
    U7 <= U148_in;
    U8 <= U149_in;
    U9 <= U150_in;

    X <= X133_in;

    Y1 <= Y116_in;
    Y2 <= Y117_in;
    Y3 <= Y118_in;
    Y4 <= Y132_in;
    Y5 <= Y133_in;
    Y6 <= Y134_in;
    Y7 <= Y148_in;
    Y8 <= Y149_in;
    Y9 <= Y150_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10000101) begin // 134

    Y133_next <= Y_onebyoneout;
    X133_next <= X_onebyoneout;

    U1 <= U117_in;
    U2 <= U118_in;
    U3 <= U119_in;
    U4 <= U133_in;
    U5 <= U134_in;
    U6 <= U135_in;
    U7 <= U149_in;
    U8 <= U150_in;
    U9 <= U151_in;

    X <= X134_in;

    Y1 <= Y117_in;
    Y2 <= Y118_in;
    Y3 <= Y119_in;
    Y4 <= Y133_in;
    Y5 <= Y134_in;
    Y6 <= Y135_in;
    Y7 <= Y149_in;
    Y8 <= Y150_in;
    Y9 <= Y151_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10000110) begin // 135

    Y134_next <= Y_onebyoneout;
    X134_next <= X_onebyoneout;

    U1 <= U118_in;
    U2 <= U119_in;
    U3 <= U120_in;
    U4 <= U134_in;
    U5 <= U135_in;
    U6 <= U136_in;
    U7 <= U150_in;
    U8 <= U151_in;
    U9 <= U152_in;

    X <= X135_in;

    Y1 <= Y118_in;
    Y2 <= Y119_in;
    Y3 <= Y120_in;
    Y4 <= Y134_in;
    Y5 <= Y135_in;
    Y6 <= Y136_in;
    Y7 <= Y150_in;
    Y8 <= Y151_in;
    Y9 <= Y152_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10000111) begin // 136

    Y135_next <= Y_onebyoneout;
    X135_next <= X_onebyoneout;

    U1 <= U119_in;
    U2 <= U120_in;
    U3 <= U121_in;
    U4 <= U135_in;
    U5 <= U136_in;
    U6 <= U137_in;
    U7 <= U151_in;
    U8 <= U152_in;
    U9 <= U153_in;

    X <= X136_in;

    Y1 <= Y119_in;
    Y2 <= Y120_in;
    Y3 <= Y121_in;
    Y4 <= Y135_in;
    Y5 <= Y136_in;
    Y6 <= Y137_in;
    Y7 <= Y151_in;
    Y8 <= Y152_in;
    Y9 <= Y153_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10001000) begin // 137

    Y136_next <= Y_onebyoneout;
    X136_next <= X_onebyoneout;

    U1 <= U120_in;
    U2 <= U121_in;
    U3 <= U122_in;
    U4 <= U136_in;
    U5 <= U137_in;
    U6 <= U138_in;
    U7 <= U152_in;
    U8 <= U153_in;
    U9 <= U154_in;

    X <= X137_in;

    Y1 <= Y120_in;
    Y2 <= Y121_in;
    Y3 <= Y122_in;
    Y4 <= Y136_in;
    Y5 <= Y137_in;
    Y6 <= Y138_in;
    Y7 <= Y152_in;
    Y8 <= Y153_in;
    Y9 <= Y154_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10001001) begin // 138

    Y137_next <= Y_onebyoneout;
    X137_next <= X_onebyoneout;

    U1 <= U121_in;
    U2 <= U122_in;
    U3 <= U123_in;
    U4 <= U137_in;
    U5 <= U138_in;
    U6 <= U139_in;
    U7 <= U153_in;
    U8 <= U154_in;
    U9 <= U155_in;

    X <= X138_in;

    Y1 <= Y121_in;
    Y2 <= Y122_in;
    Y3 <= Y123_in;
    Y4 <= Y137_in;
    Y5 <= Y138_in;
    Y6 <= Y139_in;
    Y7 <= Y153_in;
    Y8 <= Y154_in;
    Y9 <= Y155_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10001010) begin // 139

    Y138_next <= Y_onebyoneout;
    X138_next <= X_onebyoneout;

    U1 <= U122_in;
    U2 <= U123_in;
    U3 <= U124_in;
    U4 <= U138_in;
    U5 <= U139_in;
    U6 <= U140_in;
    U7 <= U154_in;
    U8 <= U155_in;
    U9 <= U156_in;

    X <= X139_in;

    Y1 <= Y122_in;
    Y2 <= Y123_in;
    Y3 <= Y124_in;
    Y4 <= Y138_in;
    Y5 <= Y139_in;
    Y6 <= Y140_in;
    Y7 <= Y154_in;
    Y8 <= Y155_in;
    Y9 <= Y156_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10001011) begin // 140

    Y139_next <= Y_onebyoneout;
    X139_next <= X_onebyoneout;

    U1 <= U123_in;
    U2 <= U124_in;
    U3 <= U125_in;
    U4 <= U139_in;
    U5 <= U140_in;
    U6 <= U141_in;
    U7 <= U155_in;
    U8 <= U156_in;
    U9 <= U157_in;

    X <= X140_in;

    Y1 <= Y123_in;
    Y2 <= Y124_in;
    Y3 <= Y125_in;
    Y4 <= Y139_in;
    Y5 <= Y140_in;
    Y6 <= Y141_in;
    Y7 <= Y155_in;
    Y8 <= Y156_in;
    Y9 <= Y157_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10001100) begin // 141

    Y140_next <= Y_onebyoneout;
    X140_next <= X_onebyoneout;

    U1 <= U124_in;
    U2 <= U125_in;
    U3 <= U126_in;
    U4 <= U140_in;
    U5 <= U141_in;
    U6 <= U142_in;
    U7 <= U156_in;
    U8 <= U157_in;
    U9 <= U158_in;

    X <= X141_in;

    Y1 <= Y124_in;
    Y2 <= Y125_in;
    Y3 <= Y126_in;
    Y4 <= Y140_in;
    Y5 <= Y141_in;
    Y6 <= Y142_in;
    Y7 <= Y156_in;
    Y8 <= Y157_in;
    Y9 <= Y158_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10001101) begin // 142

    Y141_next <= Y_onebyoneout;
    X141_next <= X_onebyoneout;

    U1 <= U125_in;
    U2 <= U126_in;
    U3 <= U127_in;
    U4 <= U141_in;
    U5 <= U142_in;
    U6 <= U143_in;
    U7 <= U157_in;
    U8 <= U158_in;
    U9 <= U159_in;

    X <= X142_in;

    Y1 <= Y125_in;
    Y2 <= Y126_in;
    Y3 <= Y127_in;
    Y4 <= Y141_in;
    Y5 <= Y142_in;
    Y6 <= Y143_in;
    Y7 <= Y157_in;
    Y8 <= Y158_in;
    Y9 <= Y159_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10001110) begin // 143

    Y142_next <= Y_onebyoneout;
    X142_next <= X_onebyoneout;

    U1 <= U126_in;
    U2 <= U127_in;
    U3 <= U128_in;
    U4 <= U142_in;
    U5 <= U143_in;
    U6 <= U144_in;
    U7 <= U158_in;
    U8 <= U159_in;
    U9 <= U160_in;

    X <= X143_in;

    Y1 <= Y126_in;
    Y2 <= Y127_in;
    Y3 <= Y128_in;
    Y4 <= Y142_in;
    Y5 <= Y143_in;
    Y6 <= Y144_in;
    Y7 <= Y158_in;
    Y8 <= Y159_in;
    Y9 <= Y160_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10001111) begin // 144

    Y143_next <= Y_onebyoneout;
    X143_next <= X_onebyoneout;

    U1 <= U127_in;
    U2 <= U128_in;
    U3 <= `WIDTH'b0;
    U4 <= U143_in;
    U5 <= U144_in;
    U6 <= `WIDTH'b0;
    U7 <= U159_in;
    U8 <= U160_in;
    U9 <= `WIDTH'b0;

    X <= X144_in;

    Y1 <= Y127_in;
    Y2 <= Y128_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y143_in;
    Y5 <= Y144_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y159_in;
    Y8 <= Y160_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10010000) begin // 145

    Y144_next <= Y_onebyoneout;
    X144_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U129_in;
    U3 <= U130_in;
    U4 <= `WIDTH'b0;
    U5 <= U145_in;
    U6 <= U146_in;
    U7 <= `WIDTH'b0;
    U8 <= U161_in;
    U9 <= U162_in;

    X <= X145_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y129_in;
    Y3 <= Y130_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y145_in;
    Y6 <= Y146_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y161_in;
    Y9 <= Y162_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10010001) begin // 146

    Y145_next <= Y_onebyoneout;
    X145_next <= X_onebyoneout;

    U1 <= U129_in;
    U2 <= U130_in;
    U3 <= U131_in;
    U4 <= U145_in;
    U5 <= U146_in;
    U6 <= U147_in;
    U7 <= U161_in;
    U8 <= U162_in;
    U9 <= U163_in;

    X <= X146_in;

    Y1 <= Y129_in;
    Y2 <= Y130_in;
    Y3 <= Y131_in;
    Y4 <= Y145_in;
    Y5 <= Y146_in;
    Y6 <= Y147_in;
    Y7 <= Y161_in;
    Y8 <= Y162_in;
    Y9 <= Y163_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10010010) begin // 147

    Y146_next <= Y_onebyoneout;
    X146_next <= X_onebyoneout;

    U1 <= U130_in;
    U2 <= U131_in;
    U3 <= U132_in;
    U4 <= U146_in;
    U5 <= U147_in;
    U6 <= U148_in;
    U7 <= U162_in;
    U8 <= U163_in;
    U9 <= U164_in;

    X <= X147_in;

    Y1 <= Y130_in;
    Y2 <= Y131_in;
    Y3 <= Y132_in;
    Y4 <= Y146_in;
    Y5 <= Y147_in;
    Y6 <= Y148_in;
    Y7 <= Y162_in;
    Y8 <= Y163_in;
    Y9 <= Y164_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10010011) begin // 148

    Y147_next <= Y_onebyoneout;
    X147_next <= X_onebyoneout;

    U1 <= U131_in;
    U2 <= U132_in;
    U3 <= U133_in;
    U4 <= U147_in;
    U5 <= U148_in;
    U6 <= U149_in;
    U7 <= U163_in;
    U8 <= U164_in;
    U9 <= U165_in;

    X <= X148_in;

    Y1 <= Y131_in;
    Y2 <= Y132_in;
    Y3 <= Y133_in;
    Y4 <= Y147_in;
    Y5 <= Y148_in;
    Y6 <= Y149_in;
    Y7 <= Y163_in;
    Y8 <= Y164_in;
    Y9 <= Y165_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10010100) begin // 149

    Y148_next <= Y_onebyoneout;
    X148_next <= X_onebyoneout;

    U1 <= U132_in;
    U2 <= U133_in;
    U3 <= U134_in;
    U4 <= U148_in;
    U5 <= U149_in;
    U6 <= U150_in;
    U7 <= U164_in;
    U8 <= U165_in;
    U9 <= U166_in;

    X <= X149_in;

    Y1 <= Y132_in;
    Y2 <= Y133_in;
    Y3 <= Y134_in;
    Y4 <= Y148_in;
    Y5 <= Y149_in;
    Y6 <= Y150_in;
    Y7 <= Y164_in;
    Y8 <= Y165_in;
    Y9 <= Y166_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10010101) begin // 150

    Y149_next <= Y_onebyoneout;
    X149_next <= X_onebyoneout;

    U1 <= U133_in;
    U2 <= U134_in;
    U3 <= U135_in;
    U4 <= U149_in;
    U5 <= U150_in;
    U6 <= U151_in;
    U7 <= U165_in;
    U8 <= U166_in;
    U9 <= U167_in;

    X <= X150_in;

    Y1 <= Y133_in;
    Y2 <= Y134_in;
    Y3 <= Y135_in;
    Y4 <= Y149_in;
    Y5 <= Y150_in;
    Y6 <= Y151_in;
    Y7 <= Y165_in;
    Y8 <= Y166_in;
    Y9 <= Y167_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10010110) begin // 151

    Y150_next <= Y_onebyoneout;
    X150_next <= X_onebyoneout;

    U1 <= U134_in;
    U2 <= U135_in;
    U3 <= U136_in;
    U4 <= U150_in;
    U5 <= U151_in;
    U6 <= U152_in;
    U7 <= U166_in;
    U8 <= U167_in;
    U9 <= U168_in;

    X <= X151_in;

    Y1 <= Y134_in;
    Y2 <= Y135_in;
    Y3 <= Y136_in;
    Y4 <= Y150_in;
    Y5 <= Y151_in;
    Y6 <= Y152_in;
    Y7 <= Y166_in;
    Y8 <= Y167_in;
    Y9 <= Y168_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10010111) begin // 152

    Y151_next <= Y_onebyoneout;
    X151_next <= X_onebyoneout;

    U1 <= U135_in;
    U2 <= U136_in;
    U3 <= U137_in;
    U4 <= U151_in;
    U5 <= U152_in;
    U6 <= U153_in;
    U7 <= U167_in;
    U8 <= U168_in;
    U9 <= U169_in;

    X <= X152_in;

    Y1 <= Y135_in;
    Y2 <= Y136_in;
    Y3 <= Y137_in;
    Y4 <= Y151_in;
    Y5 <= Y152_in;
    Y6 <= Y153_in;
    Y7 <= Y167_in;
    Y8 <= Y168_in;
    Y9 <= Y169_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10011000) begin // 153

    Y152_next <= Y_onebyoneout;
    X152_next <= X_onebyoneout;

    U1 <= U136_in;
    U2 <= U137_in;
    U3 <= U138_in;
    U4 <= U152_in;
    U5 <= U153_in;
    U6 <= U154_in;
    U7 <= U168_in;
    U8 <= U169_in;
    U9 <= U170_in;

    X <= X153_in;

    Y1 <= Y136_in;
    Y2 <= Y137_in;
    Y3 <= Y138_in;
    Y4 <= Y152_in;
    Y5 <= Y153_in;
    Y6 <= Y154_in;
    Y7 <= Y168_in;
    Y8 <= Y169_in;
    Y9 <= Y170_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10011001) begin // 154

    Y153_next <= Y_onebyoneout;
    X153_next <= X_onebyoneout;

    U1 <= U137_in;
    U2 <= U138_in;
    U3 <= U139_in;
    U4 <= U153_in;
    U5 <= U154_in;
    U6 <= U155_in;
    U7 <= U169_in;
    U8 <= U170_in;
    U9 <= U171_in;

    X <= X154_in;

    Y1 <= Y137_in;
    Y2 <= Y138_in;
    Y3 <= Y139_in;
    Y4 <= Y153_in;
    Y5 <= Y154_in;
    Y6 <= Y155_in;
    Y7 <= Y169_in;
    Y8 <= Y170_in;
    Y9 <= Y171_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10011010) begin // 155

    Y154_next <= Y_onebyoneout;
    X154_next <= X_onebyoneout;

    U1 <= U138_in;
    U2 <= U139_in;
    U3 <= U140_in;
    U4 <= U154_in;
    U5 <= U155_in;
    U6 <= U156_in;
    U7 <= U170_in;
    U8 <= U171_in;
    U9 <= U172_in;

    X <= X155_in;

    Y1 <= Y138_in;
    Y2 <= Y139_in;
    Y3 <= Y140_in;
    Y4 <= Y154_in;
    Y5 <= Y155_in;
    Y6 <= Y156_in;
    Y7 <= Y170_in;
    Y8 <= Y171_in;
    Y9 <= Y172_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10011011) begin // 156

    Y155_next <= Y_onebyoneout;
    X155_next <= X_onebyoneout;

    U1 <= U139_in;
    U2 <= U140_in;
    U3 <= U141_in;
    U4 <= U155_in;
    U5 <= U156_in;
    U6 <= U157_in;
    U7 <= U171_in;
    U8 <= U172_in;
    U9 <= U173_in;

    X <= X156_in;

    Y1 <= Y139_in;
    Y2 <= Y140_in;
    Y3 <= Y141_in;
    Y4 <= Y155_in;
    Y5 <= Y156_in;
    Y6 <= Y157_in;
    Y7 <= Y171_in;
    Y8 <= Y172_in;
    Y9 <= Y173_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10011100) begin // 157

    Y156_next <= Y_onebyoneout;
    X156_next <= X_onebyoneout;

    U1 <= U140_in;
    U2 <= U141_in;
    U3 <= U142_in;
    U4 <= U156_in;
    U5 <= U157_in;
    U6 <= U158_in;
    U7 <= U172_in;
    U8 <= U173_in;
    U9 <= U174_in;

    X <= X157_in;

    Y1 <= Y140_in;
    Y2 <= Y141_in;
    Y3 <= Y142_in;
    Y4 <= Y156_in;
    Y5 <= Y157_in;
    Y6 <= Y158_in;
    Y7 <= Y172_in;
    Y8 <= Y173_in;
    Y9 <= Y174_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10011101) begin // 158

    Y157_next <= Y_onebyoneout;
    X157_next <= X_onebyoneout;

    U1 <= U141_in;
    U2 <= U142_in;
    U3 <= U143_in;
    U4 <= U157_in;
    U5 <= U158_in;
    U6 <= U159_in;
    U7 <= U173_in;
    U8 <= U174_in;
    U9 <= U175_in;

    X <= X158_in;

    Y1 <= Y141_in;
    Y2 <= Y142_in;
    Y3 <= Y143_in;
    Y4 <= Y157_in;
    Y5 <= Y158_in;
    Y6 <= Y159_in;
    Y7 <= Y173_in;
    Y8 <= Y174_in;
    Y9 <= Y175_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10011110) begin // 159

    Y158_next <= Y_onebyoneout;
    X158_next <= X_onebyoneout;

    U1 <= U142_in;
    U2 <= U143_in;
    U3 <= U144_in;
    U4 <= U158_in;
    U5 <= U159_in;
    U6 <= U160_in;
    U7 <= U174_in;
    U8 <= U175_in;
    U9 <= U176_in;

    X <= X159_in;

    Y1 <= Y142_in;
    Y2 <= Y143_in;
    Y3 <= Y144_in;
    Y4 <= Y158_in;
    Y5 <= Y159_in;
    Y6 <= Y160_in;
    Y7 <= Y174_in;
    Y8 <= Y175_in;
    Y9 <= Y176_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10011111) begin // 160

    Y159_next <= Y_onebyoneout;
    X159_next <= X_onebyoneout;

    U1 <= U143_in;
    U2 <= U144_in;
    U3 <= `WIDTH'b0;
    U4 <= U159_in;
    U5 <= U160_in;
    U6 <= `WIDTH'b0;
    U7 <= U175_in;
    U8 <= U176_in;
    U9 <= `WIDTH'b0;

    X <= X160_in;

    Y1 <= Y143_in;
    Y2 <= Y144_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y159_in;
    Y5 <= Y160_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y175_in;
    Y8 <= Y176_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10100000) begin // 161

    Y160_next <= Y_onebyoneout;
    X160_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U145_in;
    U3 <= U146_in;
    U4 <= `WIDTH'b0;
    U5 <= U161_in;
    U6 <= U162_in;
    U7 <= `WIDTH'b0;
    U8 <= U177_in;
    U9 <= U178_in;

    X <= X161_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y145_in;
    Y3 <= Y146_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y161_in;
    Y6 <= Y162_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y177_in;
    Y9 <= Y178_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10100001) begin // 162

    Y161_next <= Y_onebyoneout;
    X161_next <= X_onebyoneout;

    U1 <= U145_in;
    U2 <= U146_in;
    U3 <= U147_in;
    U4 <= U161_in;
    U5 <= U162_in;
    U6 <= U163_in;
    U7 <= U177_in;
    U8 <= U178_in;
    U9 <= U179_in;

    X <= X162_in;

    Y1 <= Y145_in;
    Y2 <= Y146_in;
    Y3 <= Y147_in;
    Y4 <= Y161_in;
    Y5 <= Y162_in;
    Y6 <= Y163_in;
    Y7 <= Y177_in;
    Y8 <= Y178_in;
    Y9 <= Y179_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10100010) begin // 163

    Y162_next <= Y_onebyoneout;
    X162_next <= X_onebyoneout;

    U1 <= U146_in;
    U2 <= U147_in;
    U3 <= U148_in;
    U4 <= U162_in;
    U5 <= U163_in;
    U6 <= U164_in;
    U7 <= U178_in;
    U8 <= U179_in;
    U9 <= U180_in;

    X <= X163_in;

    Y1 <= Y146_in;
    Y2 <= Y147_in;
    Y3 <= Y148_in;
    Y4 <= Y162_in;
    Y5 <= Y163_in;
    Y6 <= Y164_in;
    Y7 <= Y178_in;
    Y8 <= Y179_in;
    Y9 <= Y180_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10100011) begin // 164

    Y163_next <= Y_onebyoneout;
    X163_next <= X_onebyoneout;

    U1 <= U147_in;
    U2 <= U148_in;
    U3 <= U149_in;
    U4 <= U163_in;
    U5 <= U164_in;
    U6 <= U165_in;
    U7 <= U179_in;
    U8 <= U180_in;
    U9 <= U181_in;

    X <= X164_in;

    Y1 <= Y147_in;
    Y2 <= Y148_in;
    Y3 <= Y149_in;
    Y4 <= Y163_in;
    Y5 <= Y164_in;
    Y6 <= Y165_in;
    Y7 <= Y179_in;
    Y8 <= Y180_in;
    Y9 <= Y181_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10100100) begin // 165

    Y164_next <= Y_onebyoneout;
    X164_next <= X_onebyoneout;

    U1 <= U148_in;
    U2 <= U149_in;
    U3 <= U150_in;
    U4 <= U164_in;
    U5 <= U165_in;
    U6 <= U166_in;
    U7 <= U180_in;
    U8 <= U181_in;
    U9 <= U182_in;

    X <= X165_in;

    Y1 <= Y148_in;
    Y2 <= Y149_in;
    Y3 <= Y150_in;
    Y4 <= Y164_in;
    Y5 <= Y165_in;
    Y6 <= Y166_in;
    Y7 <= Y180_in;
    Y8 <= Y181_in;
    Y9 <= Y182_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10100101) begin // 166

    Y165_next <= Y_onebyoneout;
    X165_next <= X_onebyoneout;

    U1 <= U149_in;
    U2 <= U150_in;
    U3 <= U151_in;
    U4 <= U165_in;
    U5 <= U166_in;
    U6 <= U167_in;
    U7 <= U181_in;
    U8 <= U182_in;
    U9 <= U183_in;

    X <= X166_in;

    Y1 <= Y149_in;
    Y2 <= Y150_in;
    Y3 <= Y151_in;
    Y4 <= Y165_in;
    Y5 <= Y166_in;
    Y6 <= Y167_in;
    Y7 <= Y181_in;
    Y8 <= Y182_in;
    Y9 <= Y183_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10100110) begin // 167

    Y166_next <= Y_onebyoneout;
    X166_next <= X_onebyoneout;

    U1 <= U150_in;
    U2 <= U151_in;
    U3 <= U152_in;
    U4 <= U166_in;
    U5 <= U167_in;
    U6 <= U168_in;
    U7 <= U182_in;
    U8 <= U183_in;
    U9 <= U184_in;

    X <= X167_in;

    Y1 <= Y150_in;
    Y2 <= Y151_in;
    Y3 <= Y152_in;
    Y4 <= Y166_in;
    Y5 <= Y167_in;
    Y6 <= Y168_in;
    Y7 <= Y182_in;
    Y8 <= Y183_in;
    Y9 <= Y184_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10100111) begin // 168

    Y167_next <= Y_onebyoneout;
    X167_next <= X_onebyoneout;

    U1 <= U151_in;
    U2 <= U152_in;
    U3 <= U153_in;
    U4 <= U167_in;
    U5 <= U168_in;
    U6 <= U169_in;
    U7 <= U183_in;
    U8 <= U184_in;
    U9 <= U185_in;

    X <= X168_in;

    Y1 <= Y151_in;
    Y2 <= Y152_in;
    Y3 <= Y153_in;
    Y4 <= Y167_in;
    Y5 <= Y168_in;
    Y6 <= Y169_in;
    Y7 <= Y183_in;
    Y8 <= Y184_in;
    Y9 <= Y185_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10101000) begin // 169

    Y168_next <= Y_onebyoneout;
    X168_next <= X_onebyoneout;

    U1 <= U152_in;
    U2 <= U153_in;
    U3 <= U154_in;
    U4 <= U168_in;
    U5 <= U169_in;
    U6 <= U170_in;
    U7 <= U184_in;
    U8 <= U185_in;
    U9 <= U186_in;

    X <= X169_in;

    Y1 <= Y152_in;
    Y2 <= Y153_in;
    Y3 <= Y154_in;
    Y4 <= Y168_in;
    Y5 <= Y169_in;
    Y6 <= Y170_in;
    Y7 <= Y184_in;
    Y8 <= Y185_in;
    Y9 <= Y186_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10101001) begin // 170

    Y169_next <= Y_onebyoneout;
    X169_next <= X_onebyoneout;

    U1 <= U153_in;
    U2 <= U154_in;
    U3 <= U155_in;
    U4 <= U169_in;
    U5 <= U170_in;
    U6 <= U171_in;
    U7 <= U185_in;
    U8 <= U186_in;
    U9 <= U187_in;

    X <= X170_in;

    Y1 <= Y153_in;
    Y2 <= Y154_in;
    Y3 <= Y155_in;
    Y4 <= Y169_in;
    Y5 <= Y170_in;
    Y6 <= Y171_in;
    Y7 <= Y185_in;
    Y8 <= Y186_in;
    Y9 <= Y187_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10101010) begin // 171

    Y170_next <= Y_onebyoneout;
    X170_next <= X_onebyoneout;

    U1 <= U154_in;
    U2 <= U155_in;
    U3 <= U156_in;
    U4 <= U170_in;
    U5 <= U171_in;
    U6 <= U172_in;
    U7 <= U186_in;
    U8 <= U187_in;
    U9 <= U188_in;

    X <= X171_in;

    Y1 <= Y154_in;
    Y2 <= Y155_in;
    Y3 <= Y156_in;
    Y4 <= Y170_in;
    Y5 <= Y171_in;
    Y6 <= Y172_in;
    Y7 <= Y186_in;
    Y8 <= Y187_in;
    Y9 <= Y188_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10101011) begin // 172

    Y171_next <= Y_onebyoneout;
    X171_next <= X_onebyoneout;

    U1 <= U155_in;
    U2 <= U156_in;
    U3 <= U157_in;
    U4 <= U171_in;
    U5 <= U172_in;
    U6 <= U173_in;
    U7 <= U187_in;
    U8 <= U188_in;
    U9 <= U189_in;

    X <= X172_in;

    Y1 <= Y155_in;
    Y2 <= Y156_in;
    Y3 <= Y157_in;
    Y4 <= Y171_in;
    Y5 <= Y172_in;
    Y6 <= Y173_in;
    Y7 <= Y187_in;
    Y8 <= Y188_in;
    Y9 <= Y189_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10101100) begin // 173

    Y172_next <= Y_onebyoneout;
    X172_next <= X_onebyoneout;

    U1 <= U156_in;
    U2 <= U157_in;
    U3 <= U158_in;
    U4 <= U172_in;
    U5 <= U173_in;
    U6 <= U174_in;
    U7 <= U188_in;
    U8 <= U189_in;
    U9 <= U190_in;

    X <= X173_in;

    Y1 <= Y156_in;
    Y2 <= Y157_in;
    Y3 <= Y158_in;
    Y4 <= Y172_in;
    Y5 <= Y173_in;
    Y6 <= Y174_in;
    Y7 <= Y188_in;
    Y8 <= Y189_in;
    Y9 <= Y190_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10101101) begin // 174

    Y173_next <= Y_onebyoneout;
    X173_next <= X_onebyoneout;

    U1 <= U157_in;
    U2 <= U158_in;
    U3 <= U159_in;
    U4 <= U173_in;
    U5 <= U174_in;
    U6 <= U175_in;
    U7 <= U189_in;
    U8 <= U190_in;
    U9 <= U191_in;

    X <= X174_in;

    Y1 <= Y157_in;
    Y2 <= Y158_in;
    Y3 <= Y159_in;
    Y4 <= Y173_in;
    Y5 <= Y174_in;
    Y6 <= Y175_in;
    Y7 <= Y189_in;
    Y8 <= Y190_in;
    Y9 <= Y191_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10101110) begin // 175

    Y174_next <= Y_onebyoneout;
    X174_next <= X_onebyoneout;

    U1 <= U158_in;
    U2 <= U159_in;
    U3 <= U160_in;
    U4 <= U174_in;
    U5 <= U175_in;
    U6 <= U176_in;
    U7 <= U190_in;
    U8 <= U191_in;
    U9 <= U192_in;

    X <= X175_in;

    Y1 <= Y158_in;
    Y2 <= Y159_in;
    Y3 <= Y160_in;
    Y4 <= Y174_in;
    Y5 <= Y175_in;
    Y6 <= Y176_in;
    Y7 <= Y190_in;
    Y8 <= Y191_in;
    Y9 <= Y192_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10101111) begin // 176

    Y175_next <= Y_onebyoneout;
    X175_next <= X_onebyoneout;

    U1 <= U159_in;
    U2 <= U160_in;
    U3 <= `WIDTH'b0;
    U4 <= U175_in;
    U5 <= U176_in;
    U6 <= `WIDTH'b0;
    U7 <= U191_in;
    U8 <= U192_in;
    U9 <= `WIDTH'b0;

    X <= X176_in;

    Y1 <= Y159_in;
    Y2 <= Y160_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y175_in;
    Y5 <= Y176_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y191_in;
    Y8 <= Y192_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10110000) begin // 177

    Y176_next <= Y_onebyoneout;
    X176_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U161_in;
    U3 <= U162_in;
    U4 <= `WIDTH'b0;
    U5 <= U177_in;
    U6 <= U178_in;
    U7 <= `WIDTH'b0;
    U8 <= U193_in;
    U9 <= U194_in;

    X <= X177_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y161_in;
    Y3 <= Y162_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y177_in;
    Y6 <= Y178_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y193_in;
    Y9 <= Y194_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10110001) begin // 178

    Y177_next <= Y_onebyoneout;
    X177_next <= X_onebyoneout;

    U1 <= U161_in;
    U2 <= U162_in;
    U3 <= U163_in;
    U4 <= U177_in;
    U5 <= U178_in;
    U6 <= U179_in;
    U7 <= U193_in;
    U8 <= U194_in;
    U9 <= U195_in;

    X <= X178_in;

    Y1 <= Y161_in;
    Y2 <= Y162_in;
    Y3 <= Y163_in;
    Y4 <= Y177_in;
    Y5 <= Y178_in;
    Y6 <= Y179_in;
    Y7 <= Y193_in;
    Y8 <= Y194_in;
    Y9 <= Y195_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10110010) begin // 179

    Y178_next <= Y_onebyoneout;
    X178_next <= X_onebyoneout;

    U1 <= U162_in;
    U2 <= U163_in;
    U3 <= U164_in;
    U4 <= U178_in;
    U5 <= U179_in;
    U6 <= U180_in;
    U7 <= U194_in;
    U8 <= U195_in;
    U9 <= U196_in;

    X <= X179_in;

    Y1 <= Y162_in;
    Y2 <= Y163_in;
    Y3 <= Y164_in;
    Y4 <= Y178_in;
    Y5 <= Y179_in;
    Y6 <= Y180_in;
    Y7 <= Y194_in;
    Y8 <= Y195_in;
    Y9 <= Y196_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10110011) begin // 180

    Y179_next <= Y_onebyoneout;
    X179_next <= X_onebyoneout;

    U1 <= U163_in;
    U2 <= U164_in;
    U3 <= U165_in;
    U4 <= U179_in;
    U5 <= U180_in;
    U6 <= U181_in;
    U7 <= U195_in;
    U8 <= U196_in;
    U9 <= U197_in;

    X <= X180_in;

    Y1 <= Y163_in;
    Y2 <= Y164_in;
    Y3 <= Y165_in;
    Y4 <= Y179_in;
    Y5 <= Y180_in;
    Y6 <= Y181_in;
    Y7 <= Y195_in;
    Y8 <= Y196_in;
    Y9 <= Y197_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10110100) begin // 181

    Y180_next <= Y_onebyoneout;
    X180_next <= X_onebyoneout;

    U1 <= U164_in;
    U2 <= U165_in;
    U3 <= U166_in;
    U4 <= U180_in;
    U5 <= U181_in;
    U6 <= U182_in;
    U7 <= U196_in;
    U8 <= U197_in;
    U9 <= U198_in;

    X <= X181_in;

    Y1 <= Y164_in;
    Y2 <= Y165_in;
    Y3 <= Y166_in;
    Y4 <= Y180_in;
    Y5 <= Y181_in;
    Y6 <= Y182_in;
    Y7 <= Y196_in;
    Y8 <= Y197_in;
    Y9 <= Y198_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10110101) begin // 182

    Y181_next <= Y_onebyoneout;
    X181_next <= X_onebyoneout;

    U1 <= U165_in;
    U2 <= U166_in;
    U3 <= U167_in;
    U4 <= U181_in;
    U5 <= U182_in;
    U6 <= U183_in;
    U7 <= U197_in;
    U8 <= U198_in;
    U9 <= U199_in;

    X <= X182_in;

    Y1 <= Y165_in;
    Y2 <= Y166_in;
    Y3 <= Y167_in;
    Y4 <= Y181_in;
    Y5 <= Y182_in;
    Y6 <= Y183_in;
    Y7 <= Y197_in;
    Y8 <= Y198_in;
    Y9 <= Y199_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10110110) begin // 183

    Y182_next <= Y_onebyoneout;
    X182_next <= X_onebyoneout;

    U1 <= U166_in;
    U2 <= U167_in;
    U3 <= U168_in;
    U4 <= U182_in;
    U5 <= U183_in;
    U6 <= U184_in;
    U7 <= U198_in;
    U8 <= U199_in;
    U9 <= U200_in;

    X <= X183_in;

    Y1 <= Y166_in;
    Y2 <= Y167_in;
    Y3 <= Y168_in;
    Y4 <= Y182_in;
    Y5 <= Y183_in;
    Y6 <= Y184_in;
    Y7 <= Y198_in;
    Y8 <= Y199_in;
    Y9 <= Y200_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10110111) begin // 184

    Y183_next <= Y_onebyoneout;
    X183_next <= X_onebyoneout;

    U1 <= U167_in;
    U2 <= U168_in;
    U3 <= U169_in;
    U4 <= U183_in;
    U5 <= U184_in;
    U6 <= U185_in;
    U7 <= U199_in;
    U8 <= U200_in;
    U9 <= U201_in;

    X <= X184_in;

    Y1 <= Y167_in;
    Y2 <= Y168_in;
    Y3 <= Y169_in;
    Y4 <= Y183_in;
    Y5 <= Y184_in;
    Y6 <= Y185_in;
    Y7 <= Y199_in;
    Y8 <= Y200_in;
    Y9 <= Y201_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10111000) begin // 185

    Y184_next <= Y_onebyoneout;
    X184_next <= X_onebyoneout;

    U1 <= U168_in;
    U2 <= U169_in;
    U3 <= U170_in;
    U4 <= U184_in;
    U5 <= U185_in;
    U6 <= U186_in;
    U7 <= U200_in;
    U8 <= U201_in;
    U9 <= U202_in;

    X <= X185_in;

    Y1 <= Y168_in;
    Y2 <= Y169_in;
    Y3 <= Y170_in;
    Y4 <= Y184_in;
    Y5 <= Y185_in;
    Y6 <= Y186_in;
    Y7 <= Y200_in;
    Y8 <= Y201_in;
    Y9 <= Y202_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10111001) begin // 186

    Y185_next <= Y_onebyoneout;
    X185_next <= X_onebyoneout;

    U1 <= U169_in;
    U2 <= U170_in;
    U3 <= U171_in;
    U4 <= U185_in;
    U5 <= U186_in;
    U6 <= U187_in;
    U7 <= U201_in;
    U8 <= U202_in;
    U9 <= U203_in;

    X <= X186_in;

    Y1 <= Y169_in;
    Y2 <= Y170_in;
    Y3 <= Y171_in;
    Y4 <= Y185_in;
    Y5 <= Y186_in;
    Y6 <= Y187_in;
    Y7 <= Y201_in;
    Y8 <= Y202_in;
    Y9 <= Y203_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10111010) begin // 187

    Y186_next <= Y_onebyoneout;
    X186_next <= X_onebyoneout;

    U1 <= U170_in;
    U2 <= U171_in;
    U3 <= U172_in;
    U4 <= U186_in;
    U5 <= U187_in;
    U6 <= U188_in;
    U7 <= U202_in;
    U8 <= U203_in;
    U9 <= U204_in;

    X <= X187_in;

    Y1 <= Y170_in;
    Y2 <= Y171_in;
    Y3 <= Y172_in;
    Y4 <= Y186_in;
    Y5 <= Y187_in;
    Y6 <= Y188_in;
    Y7 <= Y202_in;
    Y8 <= Y203_in;
    Y9 <= Y204_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10111011) begin // 188

    Y187_next <= Y_onebyoneout;
    X187_next <= X_onebyoneout;

    U1 <= U171_in;
    U2 <= U172_in;
    U3 <= U173_in;
    U4 <= U187_in;
    U5 <= U188_in;
    U6 <= U189_in;
    U7 <= U203_in;
    U8 <= U204_in;
    U9 <= U205_in;

    X <= X188_in;

    Y1 <= Y171_in;
    Y2 <= Y172_in;
    Y3 <= Y173_in;
    Y4 <= Y187_in;
    Y5 <= Y188_in;
    Y6 <= Y189_in;
    Y7 <= Y203_in;
    Y8 <= Y204_in;
    Y9 <= Y205_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10111100) begin // 189

    Y188_next <= Y_onebyoneout;
    X188_next <= X_onebyoneout;

    U1 <= U172_in;
    U2 <= U173_in;
    U3 <= U174_in;
    U4 <= U188_in;
    U5 <= U189_in;
    U6 <= U190_in;
    U7 <= U204_in;
    U8 <= U205_in;
    U9 <= U206_in;

    X <= X189_in;

    Y1 <= Y172_in;
    Y2 <= Y173_in;
    Y3 <= Y174_in;
    Y4 <= Y188_in;
    Y5 <= Y189_in;
    Y6 <= Y190_in;
    Y7 <= Y204_in;
    Y8 <= Y205_in;
    Y9 <= Y206_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10111101) begin // 190

    Y189_next <= Y_onebyoneout;
    X189_next <= X_onebyoneout;

    U1 <= U173_in;
    U2 <= U174_in;
    U3 <= U175_in;
    U4 <= U189_in;
    U5 <= U190_in;
    U6 <= U191_in;
    U7 <= U205_in;
    U8 <= U206_in;
    U9 <= U207_in;

    X <= X190_in;

    Y1 <= Y173_in;
    Y2 <= Y174_in;
    Y3 <= Y175_in;
    Y4 <= Y189_in;
    Y5 <= Y190_in;
    Y6 <= Y191_in;
    Y7 <= Y205_in;
    Y8 <= Y206_in;
    Y9 <= Y207_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10111110) begin // 191

    Y190_next <= Y_onebyoneout;
    X190_next <= X_onebyoneout;

    U1 <= U174_in;
    U2 <= U175_in;
    U3 <= U176_in;
    U4 <= U190_in;
    U5 <= U191_in;
    U6 <= U192_in;
    U7 <= U206_in;
    U8 <= U207_in;
    U9 <= U208_in;

    X <= X191_in;

    Y1 <= Y174_in;
    Y2 <= Y175_in;
    Y3 <= Y176_in;
    Y4 <= Y190_in;
    Y5 <= Y191_in;
    Y6 <= Y192_in;
    Y7 <= Y206_in;
    Y8 <= Y207_in;
    Y9 <= Y208_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b10111111) begin // 192

    Y191_next <= Y_onebyoneout;
    X191_next <= X_onebyoneout;

    U1 <= U175_in;
    U2 <= U176_in;
    U3 <= `WIDTH'b0;
    U4 <= U191_in;
    U5 <= U192_in;
    U6 <= `WIDTH'b0;
    U7 <= U207_in;
    U8 <= U208_in;
    U9 <= `WIDTH'b0;

    X <= X192_in;

    Y1 <= Y175_in;
    Y2 <= Y176_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y191_in;
    Y5 <= Y192_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y207_in;
    Y8 <= Y208_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11000000) begin // 193

    Y192_next <= Y_onebyoneout;
    X192_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U177_in;
    U3 <= U178_in;
    U4 <= `WIDTH'b0;
    U5 <= U193_in;
    U6 <= U194_in;
    U7 <= `WIDTH'b0;
    U8 <= U209_in;
    U9 <= U210_in;

    X <= X193_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y177_in;
    Y3 <= Y178_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y193_in;
    Y6 <= Y194_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y209_in;
    Y9 <= Y210_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11000001) begin // 194

    Y193_next <= Y_onebyoneout;
    X193_next <= X_onebyoneout;

    U1 <= U177_in;
    U2 <= U178_in;
    U3 <= U179_in;
    U4 <= U193_in;
    U5 <= U194_in;
    U6 <= U195_in;
    U7 <= U209_in;
    U8 <= U210_in;
    U9 <= U211_in;

    X <= X194_in;

    Y1 <= Y177_in;
    Y2 <= Y178_in;
    Y3 <= Y179_in;
    Y4 <= Y193_in;
    Y5 <= Y194_in;
    Y6 <= Y195_in;
    Y7 <= Y209_in;
    Y8 <= Y210_in;
    Y9 <= Y211_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11000010) begin // 195

    Y194_next <= Y_onebyoneout;
    X194_next <= X_onebyoneout;

    U1 <= U178_in;
    U2 <= U179_in;
    U3 <= U180_in;
    U4 <= U194_in;
    U5 <= U195_in;
    U6 <= U196_in;
    U7 <= U210_in;
    U8 <= U211_in;
    U9 <= U212_in;

    X <= X195_in;

    Y1 <= Y178_in;
    Y2 <= Y179_in;
    Y3 <= Y180_in;
    Y4 <= Y194_in;
    Y5 <= Y195_in;
    Y6 <= Y196_in;
    Y7 <= Y210_in;
    Y8 <= Y211_in;
    Y9 <= Y212_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11000011) begin // 196

    Y195_next <= Y_onebyoneout;
    X195_next <= X_onebyoneout;

    U1 <= U179_in;
    U2 <= U180_in;
    U3 <= U181_in;
    U4 <= U195_in;
    U5 <= U196_in;
    U6 <= U197_in;
    U7 <= U211_in;
    U8 <= U212_in;
    U9 <= U213_in;

    X <= X196_in;

    Y1 <= Y179_in;
    Y2 <= Y180_in;
    Y3 <= Y181_in;
    Y4 <= Y195_in;
    Y5 <= Y196_in;
    Y6 <= Y197_in;
    Y7 <= Y211_in;
    Y8 <= Y212_in;
    Y9 <= Y213_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11000100) begin // 197

    Y196_next <= Y_onebyoneout;
    X196_next <= X_onebyoneout;

    U1 <= U180_in;
    U2 <= U181_in;
    U3 <= U182_in;
    U4 <= U196_in;
    U5 <= U197_in;
    U6 <= U198_in;
    U7 <= U212_in;
    U8 <= U213_in;
    U9 <= U214_in;

    X <= X197_in;

    Y1 <= Y180_in;
    Y2 <= Y181_in;
    Y3 <= Y182_in;
    Y4 <= Y196_in;
    Y5 <= Y197_in;
    Y6 <= Y198_in;
    Y7 <= Y212_in;
    Y8 <= Y213_in;
    Y9 <= Y214_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11000101) begin // 198

    Y197_next <= Y_onebyoneout;
    X197_next <= X_onebyoneout;

    U1 <= U181_in;
    U2 <= U182_in;
    U3 <= U183_in;
    U4 <= U197_in;
    U5 <= U198_in;
    U6 <= U199_in;
    U7 <= U213_in;
    U8 <= U214_in;
    U9 <= U215_in;

    X <= X198_in;

    Y1 <= Y181_in;
    Y2 <= Y182_in;
    Y3 <= Y183_in;
    Y4 <= Y197_in;
    Y5 <= Y198_in;
    Y6 <= Y199_in;
    Y7 <= Y213_in;
    Y8 <= Y214_in;
    Y9 <= Y215_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11000110) begin // 199

    Y198_next <= Y_onebyoneout;
    X198_next <= X_onebyoneout;

    U1 <= U182_in;
    U2 <= U183_in;
    U3 <= U184_in;
    U4 <= U198_in;
    U5 <= U199_in;
    U6 <= U200_in;
    U7 <= U214_in;
    U8 <= U215_in;
    U9 <= U216_in;

    X <= X199_in;

    Y1 <= Y182_in;
    Y2 <= Y183_in;
    Y3 <= Y184_in;
    Y4 <= Y198_in;
    Y5 <= Y199_in;
    Y6 <= Y200_in;
    Y7 <= Y214_in;
    Y8 <= Y215_in;
    Y9 <= Y216_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11000111) begin // 200

    Y199_next <= Y_onebyoneout;
    X199_next <= X_onebyoneout;

    U1 <= U183_in;
    U2 <= U184_in;
    U3 <= U185_in;
    U4 <= U199_in;
    U5 <= U200_in;
    U6 <= U201_in;
    U7 <= U215_in;
    U8 <= U216_in;
    U9 <= U217_in;

    X <= X200_in;

    Y1 <= Y183_in;
    Y2 <= Y184_in;
    Y3 <= Y185_in;
    Y4 <= Y199_in;
    Y5 <= Y200_in;
    Y6 <= Y201_in;
    Y7 <= Y215_in;
    Y8 <= Y216_in;
    Y9 <= Y217_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11001000) begin // 201

    Y200_next <= Y_onebyoneout;
    X200_next <= X_onebyoneout;

    U1 <= U184_in;
    U2 <= U185_in;
    U3 <= U186_in;
    U4 <= U200_in;
    U5 <= U201_in;
    U6 <= U202_in;
    U7 <= U216_in;
    U8 <= U217_in;
    U9 <= U218_in;

    X <= X201_in;

    Y1 <= Y184_in;
    Y2 <= Y185_in;
    Y3 <= Y186_in;
    Y4 <= Y200_in;
    Y5 <= Y201_in;
    Y6 <= Y202_in;
    Y7 <= Y216_in;
    Y8 <= Y217_in;
    Y9 <= Y218_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11001001) begin // 202

    Y201_next <= Y_onebyoneout;
    X201_next <= X_onebyoneout;

    U1 <= U185_in;
    U2 <= U186_in;
    U3 <= U187_in;
    U4 <= U201_in;
    U5 <= U202_in;
    U6 <= U203_in;
    U7 <= U217_in;
    U8 <= U218_in;
    U9 <= U219_in;

    X <= X202_in;

    Y1 <= Y185_in;
    Y2 <= Y186_in;
    Y3 <= Y187_in;
    Y4 <= Y201_in;
    Y5 <= Y202_in;
    Y6 <= Y203_in;
    Y7 <= Y217_in;
    Y8 <= Y218_in;
    Y9 <= Y219_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11001010) begin // 203

    Y202_next <= Y_onebyoneout;
    X202_next <= X_onebyoneout;

    U1 <= U186_in;
    U2 <= U187_in;
    U3 <= U188_in;
    U4 <= U202_in;
    U5 <= U203_in;
    U6 <= U204_in;
    U7 <= U218_in;
    U8 <= U219_in;
    U9 <= U220_in;

    X <= X203_in;

    Y1 <= Y186_in;
    Y2 <= Y187_in;
    Y3 <= Y188_in;
    Y4 <= Y202_in;
    Y5 <= Y203_in;
    Y6 <= Y204_in;
    Y7 <= Y218_in;
    Y8 <= Y219_in;
    Y9 <= Y220_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11001011) begin // 204

    Y203_next <= Y_onebyoneout;
    X203_next <= X_onebyoneout;

    U1 <= U187_in;
    U2 <= U188_in;
    U3 <= U189_in;
    U4 <= U203_in;
    U5 <= U204_in;
    U6 <= U205_in;
    U7 <= U219_in;
    U8 <= U220_in;
    U9 <= U221_in;

    X <= X204_in;

    Y1 <= Y187_in;
    Y2 <= Y188_in;
    Y3 <= Y189_in;
    Y4 <= Y203_in;
    Y5 <= Y204_in;
    Y6 <= Y205_in;
    Y7 <= Y219_in;
    Y8 <= Y220_in;
    Y9 <= Y221_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11001100) begin // 205

    Y204_next <= Y_onebyoneout;
    X204_next <= X_onebyoneout;

    U1 <= U188_in;
    U2 <= U189_in;
    U3 <= U190_in;
    U4 <= U204_in;
    U5 <= U205_in;
    U6 <= U206_in;
    U7 <= U220_in;
    U8 <= U221_in;
    U9 <= U222_in;

    X <= X205_in;

    Y1 <= Y188_in;
    Y2 <= Y189_in;
    Y3 <= Y190_in;
    Y4 <= Y204_in;
    Y5 <= Y205_in;
    Y6 <= Y206_in;
    Y7 <= Y220_in;
    Y8 <= Y221_in;
    Y9 <= Y222_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11001101) begin // 206

    Y205_next <= Y_onebyoneout;
    X205_next <= X_onebyoneout;

    U1 <= U189_in;
    U2 <= U190_in;
    U3 <= U191_in;
    U4 <= U205_in;
    U5 <= U206_in;
    U6 <= U207_in;
    U7 <= U221_in;
    U8 <= U222_in;
    U9 <= U223_in;

    X <= X206_in;

    Y1 <= Y189_in;
    Y2 <= Y190_in;
    Y3 <= Y191_in;
    Y4 <= Y205_in;
    Y5 <= Y206_in;
    Y6 <= Y207_in;
    Y7 <= Y221_in;
    Y8 <= Y222_in;
    Y9 <= Y223_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11001110) begin // 207

    Y206_next <= Y_onebyoneout;
    X206_next <= X_onebyoneout;

    U1 <= U190_in;
    U2 <= U191_in;
    U3 <= U192_in;
    U4 <= U206_in;
    U5 <= U207_in;
    U6 <= U208_in;
    U7 <= U222_in;
    U8 <= U223_in;
    U9 <= U224_in;

    X <= X207_in;

    Y1 <= Y190_in;
    Y2 <= Y191_in;
    Y3 <= Y192_in;
    Y4 <= Y206_in;
    Y5 <= Y207_in;
    Y6 <= Y208_in;
    Y7 <= Y222_in;
    Y8 <= Y223_in;
    Y9 <= Y224_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11001111) begin // 208

    Y207_next <= Y_onebyoneout;
    X207_next <= X_onebyoneout;

    U1 <= U191_in;
    U2 <= U192_in;
    U3 <= `WIDTH'b0;
    U4 <= U207_in;
    U5 <= U208_in;
    U6 <= `WIDTH'b0;
    U7 <= U223_in;
    U8 <= U224_in;
    U9 <= `WIDTH'b0;

    X <= X208_in;

    Y1 <= Y191_in;
    Y2 <= Y192_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y207_in;
    Y5 <= Y208_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y223_in;
    Y8 <= Y224_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11010000) begin // 209

    Y208_next <= Y_onebyoneout;
    X208_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U193_in;
    U3 <= U194_in;
    U4 <= `WIDTH'b0;
    U5 <= U209_in;
    U6 <= U210_in;
    U7 <= `WIDTH'b0;
    U8 <= U225_in;
    U9 <= U226_in;

    X <= X209_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y193_in;
    Y3 <= Y194_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y209_in;
    Y6 <= Y210_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y225_in;
    Y9 <= Y226_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11010001) begin // 210

    Y209_next <= Y_onebyoneout;
    X209_next <= X_onebyoneout;

    U1 <= U193_in;
    U2 <= U194_in;
    U3 <= U195_in;
    U4 <= U209_in;
    U5 <= U210_in;
    U6 <= U211_in;
    U7 <= U225_in;
    U8 <= U226_in;
    U9 <= U227_in;

    X <= X210_in;

    Y1 <= Y193_in;
    Y2 <= Y194_in;
    Y3 <= Y195_in;
    Y4 <= Y209_in;
    Y5 <= Y210_in;
    Y6 <= Y211_in;
    Y7 <= Y225_in;
    Y8 <= Y226_in;
    Y9 <= Y227_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11010010) begin // 211

    Y210_next <= Y_onebyoneout;
    X210_next <= X_onebyoneout;

    U1 <= U194_in;
    U2 <= U195_in;
    U3 <= U196_in;
    U4 <= U210_in;
    U5 <= U211_in;
    U6 <= U212_in;
    U7 <= U226_in;
    U8 <= U227_in;
    U9 <= U228_in;

    X <= X211_in;

    Y1 <= Y194_in;
    Y2 <= Y195_in;
    Y3 <= Y196_in;
    Y4 <= Y210_in;
    Y5 <= Y211_in;
    Y6 <= Y212_in;
    Y7 <= Y226_in;
    Y8 <= Y227_in;
    Y9 <= Y228_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11010011) begin // 212

    Y211_next <= Y_onebyoneout;
    X211_next <= X_onebyoneout;

    U1 <= U195_in;
    U2 <= U196_in;
    U3 <= U197_in;
    U4 <= U211_in;
    U5 <= U212_in;
    U6 <= U213_in;
    U7 <= U227_in;
    U8 <= U228_in;
    U9 <= U229_in;

    X <= X212_in;

    Y1 <= Y195_in;
    Y2 <= Y196_in;
    Y3 <= Y197_in;
    Y4 <= Y211_in;
    Y5 <= Y212_in;
    Y6 <= Y213_in;
    Y7 <= Y227_in;
    Y8 <= Y228_in;
    Y9 <= Y229_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11010100) begin // 213

    Y212_next <= Y_onebyoneout;
    X212_next <= X_onebyoneout;

    U1 <= U196_in;
    U2 <= U197_in;
    U3 <= U198_in;
    U4 <= U212_in;
    U5 <= U213_in;
    U6 <= U214_in;
    U7 <= U228_in;
    U8 <= U229_in;
    U9 <= U230_in;

    X <= X213_in;

    Y1 <= Y196_in;
    Y2 <= Y197_in;
    Y3 <= Y198_in;
    Y4 <= Y212_in;
    Y5 <= Y213_in;
    Y6 <= Y214_in;
    Y7 <= Y228_in;
    Y8 <= Y229_in;
    Y9 <= Y230_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11010101) begin // 214

    Y213_next <= Y_onebyoneout;
    X213_next <= X_onebyoneout;

    U1 <= U197_in;
    U2 <= U198_in;
    U3 <= U199_in;
    U4 <= U213_in;
    U5 <= U214_in;
    U6 <= U215_in;
    U7 <= U229_in;
    U8 <= U230_in;
    U9 <= U231_in;

    X <= X214_in;

    Y1 <= Y197_in;
    Y2 <= Y198_in;
    Y3 <= Y199_in;
    Y4 <= Y213_in;
    Y5 <= Y214_in;
    Y6 <= Y215_in;
    Y7 <= Y229_in;
    Y8 <= Y230_in;
    Y9 <= Y231_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11010110) begin // 215

    Y214_next <= Y_onebyoneout;
    X214_next <= X_onebyoneout;

    U1 <= U198_in;
    U2 <= U199_in;
    U3 <= U200_in;
    U4 <= U214_in;
    U5 <= U215_in;
    U6 <= U216_in;
    U7 <= U230_in;
    U8 <= U231_in;
    U9 <= U232_in;

    X <= X215_in;

    Y1 <= Y198_in;
    Y2 <= Y199_in;
    Y3 <= Y200_in;
    Y4 <= Y214_in;
    Y5 <= Y215_in;
    Y6 <= Y216_in;
    Y7 <= Y230_in;
    Y8 <= Y231_in;
    Y9 <= Y232_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11010111) begin // 216

    Y215_next <= Y_onebyoneout;
    X215_next <= X_onebyoneout;

    U1 <= U199_in;
    U2 <= U200_in;
    U3 <= U201_in;
    U4 <= U215_in;
    U5 <= U216_in;
    U6 <= U217_in;
    U7 <= U231_in;
    U8 <= U232_in;
    U9 <= U233_in;

    X <= X216_in;

    Y1 <= Y199_in;
    Y2 <= Y200_in;
    Y3 <= Y201_in;
    Y4 <= Y215_in;
    Y5 <= Y216_in;
    Y6 <= Y217_in;
    Y7 <= Y231_in;
    Y8 <= Y232_in;
    Y9 <= Y233_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11011000) begin // 217

    Y216_next <= Y_onebyoneout;
    X216_next <= X_onebyoneout;

    U1 <= U200_in;
    U2 <= U201_in;
    U3 <= U202_in;
    U4 <= U216_in;
    U5 <= U217_in;
    U6 <= U218_in;
    U7 <= U232_in;
    U8 <= U233_in;
    U9 <= U234_in;

    X <= X217_in;

    Y1 <= Y200_in;
    Y2 <= Y201_in;
    Y3 <= Y202_in;
    Y4 <= Y216_in;
    Y5 <= Y217_in;
    Y6 <= Y218_in;
    Y7 <= Y232_in;
    Y8 <= Y233_in;
    Y9 <= Y234_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11011001) begin // 218

    Y217_next <= Y_onebyoneout;
    X217_next <= X_onebyoneout;

    U1 <= U201_in;
    U2 <= U202_in;
    U3 <= U203_in;
    U4 <= U217_in;
    U5 <= U218_in;
    U6 <= U219_in;
    U7 <= U233_in;
    U8 <= U234_in;
    U9 <= U235_in;

    X <= X218_in;

    Y1 <= Y201_in;
    Y2 <= Y202_in;
    Y3 <= Y203_in;
    Y4 <= Y217_in;
    Y5 <= Y218_in;
    Y6 <= Y219_in;
    Y7 <= Y233_in;
    Y8 <= Y234_in;
    Y9 <= Y235_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11011010) begin // 219

    Y218_next <= Y_onebyoneout;
    X218_next <= X_onebyoneout;

    U1 <= U202_in;
    U2 <= U203_in;
    U3 <= U204_in;
    U4 <= U218_in;
    U5 <= U219_in;
    U6 <= U220_in;
    U7 <= U234_in;
    U8 <= U235_in;
    U9 <= U236_in;

    X <= X219_in;

    Y1 <= Y202_in;
    Y2 <= Y203_in;
    Y3 <= Y204_in;
    Y4 <= Y218_in;
    Y5 <= Y219_in;
    Y6 <= Y220_in;
    Y7 <= Y234_in;
    Y8 <= Y235_in;
    Y9 <= Y236_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11011011) begin // 220

    Y219_next <= Y_onebyoneout;
    X219_next <= X_onebyoneout;

    U1 <= U203_in;
    U2 <= U204_in;
    U3 <= U205_in;
    U4 <= U219_in;
    U5 <= U220_in;
    U6 <= U221_in;
    U7 <= U235_in;
    U8 <= U236_in;
    U9 <= U237_in;

    X <= X220_in;

    Y1 <= Y203_in;
    Y2 <= Y204_in;
    Y3 <= Y205_in;
    Y4 <= Y219_in;
    Y5 <= Y220_in;
    Y6 <= Y221_in;
    Y7 <= Y235_in;
    Y8 <= Y236_in;
    Y9 <= Y237_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11011100) begin // 221

    Y220_next <= Y_onebyoneout;
    X220_next <= X_onebyoneout;

    U1 <= U204_in;
    U2 <= U205_in;
    U3 <= U206_in;
    U4 <= U220_in;
    U5 <= U221_in;
    U6 <= U222_in;
    U7 <= U236_in;
    U8 <= U237_in;
    U9 <= U238_in;

    X <= X221_in;

    Y1 <= Y204_in;
    Y2 <= Y205_in;
    Y3 <= Y206_in;
    Y4 <= Y220_in;
    Y5 <= Y221_in;
    Y6 <= Y222_in;
    Y7 <= Y236_in;
    Y8 <= Y237_in;
    Y9 <= Y238_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11011101) begin // 222

    Y221_next <= Y_onebyoneout;
    X221_next <= X_onebyoneout;

    U1 <= U205_in;
    U2 <= U206_in;
    U3 <= U207_in;
    U4 <= U221_in;
    U5 <= U222_in;
    U6 <= U223_in;
    U7 <= U237_in;
    U8 <= U238_in;
    U9 <= U239_in;

    X <= X222_in;

    Y1 <= Y205_in;
    Y2 <= Y206_in;
    Y3 <= Y207_in;
    Y4 <= Y221_in;
    Y5 <= Y222_in;
    Y6 <= Y223_in;
    Y7 <= Y237_in;
    Y8 <= Y238_in;
    Y9 <= Y239_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11011110) begin // 223

    Y222_next <= Y_onebyoneout;
    X222_next <= X_onebyoneout;

    U1 <= U206_in;
    U2 <= U207_in;
    U3 <= U208_in;
    U4 <= U222_in;
    U5 <= U223_in;
    U6 <= U224_in;
    U7 <= U238_in;
    U8 <= U239_in;
    U9 <= U240_in;

    X <= X223_in;

    Y1 <= Y206_in;
    Y2 <= Y207_in;
    Y3 <= Y208_in;
    Y4 <= Y222_in;
    Y5 <= Y223_in;
    Y6 <= Y224_in;
    Y7 <= Y238_in;
    Y8 <= Y239_in;
    Y9 <= Y240_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11011111) begin // 224

    Y223_next <= Y_onebyoneout;
    X223_next <= X_onebyoneout;

    U1 <= U207_in;
    U2 <= U208_in;
    U3 <= `WIDTH'b0;
    U4 <= U223_in;
    U5 <= U224_in;
    U6 <= `WIDTH'b0;
    U7 <= U239_in;
    U8 <= U240_in;
    U9 <= `WIDTH'b0;

    X <= X224_in;

    Y1 <= Y207_in;
    Y2 <= Y208_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y223_in;
    Y5 <= Y224_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y239_in;
    Y8 <= Y240_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11100000) begin // 225

    Y224_next <= Y_onebyoneout;
    X224_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U209_in;
    U3 <= U210_in;
    U4 <= `WIDTH'b0;
    U5 <= U225_in;
    U6 <= U226_in;
    U7 <= `WIDTH'b0;
    U8 <= U241_in;
    U9 <= U242_in;

    X <= X225_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y209_in;
    Y3 <= Y210_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y225_in;
    Y6 <= Y226_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= Y241_in;
    Y9 <= Y242_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11100001) begin // 226

    Y225_next <= Y_onebyoneout;
    X225_next <= X_onebyoneout;

    U1 <= U209_in;
    U2 <= U210_in;
    U3 <= U211_in;
    U4 <= U225_in;
    U5 <= U226_in;
    U6 <= U227_in;
    U7 <= U241_in;
    U8 <= U242_in;
    U9 <= U243_in;

    X <= X226_in;

    Y1 <= Y209_in;
    Y2 <= Y210_in;
    Y3 <= Y211_in;
    Y4 <= Y225_in;
    Y5 <= Y226_in;
    Y6 <= Y227_in;
    Y7 <= Y241_in;
    Y8 <= Y242_in;
    Y9 <= Y243_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11100010) begin // 227

    Y226_next <= Y_onebyoneout;
    X226_next <= X_onebyoneout;

    U1 <= U210_in;
    U2 <= U211_in;
    U3 <= U212_in;
    U4 <= U226_in;
    U5 <= U227_in;
    U6 <= U228_in;
    U7 <= U242_in;
    U8 <= U243_in;
    U9 <= U244_in;

    X <= X227_in;

    Y1 <= Y210_in;
    Y2 <= Y211_in;
    Y3 <= Y212_in;
    Y4 <= Y226_in;
    Y5 <= Y227_in;
    Y6 <= Y228_in;
    Y7 <= Y242_in;
    Y8 <= Y243_in;
    Y9 <= Y244_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11100011) begin // 228

    Y227_next <= Y_onebyoneout;
    X227_next <= X_onebyoneout;

    U1 <= U211_in;
    U2 <= U212_in;
    U3 <= U213_in;
    U4 <= U227_in;
    U5 <= U228_in;
    U6 <= U229_in;
    U7 <= U243_in;
    U8 <= U244_in;
    U9 <= U245_in;

    X <= X228_in;

    Y1 <= Y211_in;
    Y2 <= Y212_in;
    Y3 <= Y213_in;
    Y4 <= Y227_in;
    Y5 <= Y228_in;
    Y6 <= Y229_in;
    Y7 <= Y243_in;
    Y8 <= Y244_in;
    Y9 <= Y245_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11100100) begin // 229

    Y228_next <= Y_onebyoneout;
    X228_next <= X_onebyoneout;

    U1 <= U212_in;
    U2 <= U213_in;
    U3 <= U214_in;
    U4 <= U228_in;
    U5 <= U229_in;
    U6 <= U230_in;
    U7 <= U244_in;
    U8 <= U245_in;
    U9 <= U246_in;

    X <= X229_in;

    Y1 <= Y212_in;
    Y2 <= Y213_in;
    Y3 <= Y214_in;
    Y4 <= Y228_in;
    Y5 <= Y229_in;
    Y6 <= Y230_in;
    Y7 <= Y244_in;
    Y8 <= Y245_in;
    Y9 <= Y246_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11100101) begin // 230

    Y229_next <= Y_onebyoneout;
    X229_next <= X_onebyoneout;

    U1 <= U213_in;
    U2 <= U214_in;
    U3 <= U215_in;
    U4 <= U229_in;
    U5 <= U230_in;
    U6 <= U231_in;
    U7 <= U245_in;
    U8 <= U246_in;
    U9 <= U247_in;

    X <= X230_in;

    Y1 <= Y213_in;
    Y2 <= Y214_in;
    Y3 <= Y215_in;
    Y4 <= Y229_in;
    Y5 <= Y230_in;
    Y6 <= Y231_in;
    Y7 <= Y245_in;
    Y8 <= Y246_in;
    Y9 <= Y247_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11100110) begin // 231

    Y230_next <= Y_onebyoneout;
    X230_next <= X_onebyoneout;

    U1 <= U214_in;
    U2 <= U215_in;
    U3 <= U216_in;
    U4 <= U230_in;
    U5 <= U231_in;
    U6 <= U232_in;
    U7 <= U246_in;
    U8 <= U247_in;
    U9 <= U248_in;

    X <= X231_in;

    Y1 <= Y214_in;
    Y2 <= Y215_in;
    Y3 <= Y216_in;
    Y4 <= Y230_in;
    Y5 <= Y231_in;
    Y6 <= Y232_in;
    Y7 <= Y246_in;
    Y8 <= Y247_in;
    Y9 <= Y248_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11100111) begin // 232

    Y231_next <= Y_onebyoneout;
    X231_next <= X_onebyoneout;

    U1 <= U215_in;
    U2 <= U216_in;
    U3 <= U217_in;
    U4 <= U231_in;
    U5 <= U232_in;
    U6 <= U233_in;
    U7 <= U247_in;
    U8 <= U248_in;
    U9 <= U249_in;

    X <= X232_in;

    Y1 <= Y215_in;
    Y2 <= Y216_in;
    Y3 <= Y217_in;
    Y4 <= Y231_in;
    Y5 <= Y232_in;
    Y6 <= Y233_in;
    Y7 <= Y247_in;
    Y8 <= Y248_in;
    Y9 <= Y249_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11101000) begin // 233

    Y232_next <= Y_onebyoneout;
    X232_next <= X_onebyoneout;

    U1 <= U216_in;
    U2 <= U217_in;
    U3 <= U218_in;
    U4 <= U232_in;
    U5 <= U233_in;
    U6 <= U234_in;
    U7 <= U248_in;
    U8 <= U249_in;
    U9 <= U250_in;

    X <= X233_in;

    Y1 <= Y216_in;
    Y2 <= Y217_in;
    Y3 <= Y218_in;
    Y4 <= Y232_in;
    Y5 <= Y233_in;
    Y6 <= Y234_in;
    Y7 <= Y248_in;
    Y8 <= Y249_in;
    Y9 <= Y250_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11101001) begin // 234

    Y233_next <= Y_onebyoneout;
    X233_next <= X_onebyoneout;

    U1 <= U217_in;
    U2 <= U218_in;
    U3 <= U219_in;
    U4 <= U233_in;
    U5 <= U234_in;
    U6 <= U235_in;
    U7 <= U249_in;
    U8 <= U250_in;
    U9 <= U251_in;

    X <= X234_in;

    Y1 <= Y217_in;
    Y2 <= Y218_in;
    Y3 <= Y219_in;
    Y4 <= Y233_in;
    Y5 <= Y234_in;
    Y6 <= Y235_in;
    Y7 <= Y249_in;
    Y8 <= Y250_in;
    Y9 <= Y251_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11101010) begin // 235

    Y234_next <= Y_onebyoneout;
    X234_next <= X_onebyoneout;

    U1 <= U218_in;
    U2 <= U219_in;
    U3 <= U220_in;
    U4 <= U234_in;
    U5 <= U235_in;
    U6 <= U236_in;
    U7 <= U250_in;
    U8 <= U251_in;
    U9 <= U252_in;

    X <= X235_in;

    Y1 <= Y218_in;
    Y2 <= Y219_in;
    Y3 <= Y220_in;
    Y4 <= Y234_in;
    Y5 <= Y235_in;
    Y6 <= Y236_in;
    Y7 <= Y250_in;
    Y8 <= Y251_in;
    Y9 <= Y252_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11101011) begin // 236

    Y235_next <= Y_onebyoneout;
    X235_next <= X_onebyoneout;

    U1 <= U219_in;
    U2 <= U220_in;
    U3 <= U221_in;
    U4 <= U235_in;
    U5 <= U236_in;
    U6 <= U237_in;
    U7 <= U251_in;
    U8 <= U252_in;
    U9 <= U253_in;

    X <= X236_in;

    Y1 <= Y219_in;
    Y2 <= Y220_in;
    Y3 <= Y221_in;
    Y4 <= Y235_in;
    Y5 <= Y236_in;
    Y6 <= Y237_in;
    Y7 <= Y251_in;
    Y8 <= Y252_in;
    Y9 <= Y253_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11101100) begin // 237

    Y236_next <= Y_onebyoneout;
    X236_next <= X_onebyoneout;

    U1 <= U220_in;
    U2 <= U221_in;
    U3 <= U222_in;
    U4 <= U236_in;
    U5 <= U237_in;
    U6 <= U238_in;
    U7 <= U252_in;
    U8 <= U253_in;
    U9 <= U254_in;

    X <= X237_in;

    Y1 <= Y220_in;
    Y2 <= Y221_in;
    Y3 <= Y222_in;
    Y4 <= Y236_in;
    Y5 <= Y237_in;
    Y6 <= Y238_in;
    Y7 <= Y252_in;
    Y8 <= Y253_in;
    Y9 <= Y254_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11101101) begin // 238

    Y237_next <= Y_onebyoneout;
    X237_next <= X_onebyoneout;

    U1 <= U221_in;
    U2 <= U222_in;
    U3 <= U223_in;
    U4 <= U237_in;
    U5 <= U238_in;
    U6 <= U239_in;
    U7 <= U253_in;
    U8 <= U254_in;
    U9 <= U255_in;

    X <= X238_in;

    Y1 <= Y221_in;
    Y2 <= Y222_in;
    Y3 <= Y223_in;
    Y4 <= Y237_in;
    Y5 <= Y238_in;
    Y6 <= Y239_in;
    Y7 <= Y253_in;
    Y8 <= Y254_in;
    Y9 <= Y255_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11101110) begin // 239

    Y238_next <= Y_onebyoneout;
    X238_next <= X_onebyoneout;

    U1 <= U222_in;
    U2 <= U223_in;
    U3 <= U224_in;
    U4 <= U238_in;
    U5 <= U239_in;
    U6 <= U240_in;
    U7 <= U254_in;
    U8 <= U255_in;
    U9 <= U256_in;

    X <= X239_in;

    Y1 <= Y222_in;
    Y2 <= Y223_in;
    Y3 <= Y224_in;
    Y4 <= Y238_in;
    Y5 <= Y239_in;
    Y6 <= Y240_in;
    Y7 <= Y254_in;
    Y8 <= Y255_in;
    Y9 <= Y256_in;


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11101111) begin // 240

    Y239_next <= Y_onebyoneout;
    X239_next <= X_onebyoneout;

    U1 <= U223_in;
    U2 <= U224_in;
    U3 <= `WIDTH'b0;
    U4 <= U239_in;
    U5 <= U240_in;
    U6 <= `WIDTH'b0;
    U7 <= U255_in;
    U8 <= U256_in;
    U9 <= `WIDTH'b0;

    X <= X240_in;

    Y1 <= Y223_in;
    Y2 <= Y224_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y239_in;
    Y5 <= Y240_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= Y255_in;
    Y8 <= Y256_in;
    Y9 <= {(2 * `WIDTH){1'b0}};

  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11110000) begin // 241

    Y240_next <= Y_onebyoneout;
    X240_next <= X_onebyoneout;

    U1 <= `WIDTH'b0;
    U2 <= U225_in;
    U3 <= U226_in;
    U4 <= `WIDTH'b0;
    U5 <= U241_in;
    U6 <= U242_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X241_in;

    Y1 <= {(2 * `WIDTH){1'b0}};
    Y2 <= Y225_in;
    Y3 <= Y226_in;
    Y4 <= {(2 * `WIDTH){1'b0}};
    Y5 <= Y241_in;
    Y6 <= Y242_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11110001) begin // 242

    Y241_next <= Y_onebyoneout;
    X241_next <= X_onebyoneout;

    U1 <= U225_in;
    U2 <= U226_in;
    U3 <= U227_in;
    U4 <= U241_in;
    U5 <= U242_in;
    U6 <= U243_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X242_in;

    Y1 <= Y225_in;
    Y2 <= Y226_in;
    Y3 <= Y227_in;
    Y4 <= Y241_in;
    Y5 <= Y242_in;
    Y6 <= Y243_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11110010) begin // 243

    Y242_next <= Y_onebyoneout;
    X242_next <= X_onebyoneout;

    U1 <= U226_in;
    U2 <= U227_in;
    U3 <= U228_in;
    U4 <= U242_in;
    U5 <= U243_in;
    U6 <= U244_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X243_in;

    Y1 <= Y226_in;
    Y2 <= Y227_in;
    Y3 <= Y228_in;
    Y4 <= Y242_in;
    Y5 <= Y243_in;
    Y6 <= Y244_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11110011) begin // 244

    Y243_next <= Y_onebyoneout;
    X243_next <= X_onebyoneout;

    U1 <= U227_in;
    U2 <= U228_in;
    U3 <= U229_in;
    U4 <= U243_in;
    U5 <= U244_in;
    U6 <= U245_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X244_in;

    Y1 <= Y227_in;
    Y2 <= Y228_in;
    Y3 <= Y229_in;
    Y4 <= Y243_in;
    Y5 <= Y244_in;
    Y6 <= Y245_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11110100) begin // 245

    Y244_next <= Y_onebyoneout;
    X244_next <= X_onebyoneout;

    U1 <= U228_in;
    U2 <= U229_in;
    U3 <= U230_in;
    U4 <= U244_in;
    U5 <= U245_in;
    U6 <= U246_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X245_in;

    Y1 <= Y228_in;
    Y2 <= Y229_in;
    Y3 <= Y230_in;
    Y4 <= Y244_in;
    Y5 <= Y245_in;
    Y6 <= Y246_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11110101) begin // 246

    Y245_next <= Y_onebyoneout;
    X245_next <= X_onebyoneout;

    U1 <= U229_in;
    U2 <= U230_in;
    U3 <= U231_in;
    U4 <= U245_in;
    U5 <= U246_in;
    U6 <= U247_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X246_in;

    Y1 <= Y229_in;
    Y2 <= Y230_in;
    Y3 <= Y231_in;
    Y4 <= Y245_in;
    Y5 <= Y246_in;
    Y6 <= Y247_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11110110) begin // 247

    Y246_next <= Y_onebyoneout;
    X246_next <= X_onebyoneout;

    U1 <= U230_in;
    U2 <= U231_in;
    U3 <= U232_in;
    U4 <= U246_in;
    U5 <= U247_in;
    U6 <= U248_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X247_in;

    Y1 <= Y230_in;
    Y2 <= Y231_in;
    Y3 <= Y232_in;
    Y4 <= Y246_in;
    Y5 <= Y247_in;
    Y6 <= Y248_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11110111) begin // 248

    Y247_next <= Y_onebyoneout;
    X247_next <= X_onebyoneout;

    U1 <= U231_in;
    U2 <= U232_in;
    U3 <= U233_in;
    U4 <= U247_in;
    U5 <= U248_in;
    U6 <= U249_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X248_in;

    Y1 <= Y231_in;
    Y2 <= Y232_in;
    Y3 <= Y233_in;
    Y4 <= Y247_in;
    Y5 <= Y248_in;
    Y6 <= Y249_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11111000) begin // 249

    Y248_next <= Y_onebyoneout;
    X248_next <= X_onebyoneout;

    U1 <= U232_in;
    U2 <= U233_in;
    U3 <= U234_in;
    U4 <= U248_in;
    U5 <= U249_in;
    U6 <= U250_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X249_in;

    Y1 <= Y232_in;
    Y2 <= Y233_in;
    Y3 <= Y234_in;
    Y4 <= Y248_in;
    Y5 <= Y249_in;
    Y6 <= Y250_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11111001) begin // 250

    Y249_next <= Y_onebyoneout;
    X249_next <= X_onebyoneout;

    U1 <= U233_in;
    U2 <= U234_in;
    U3 <= U235_in;
    U4 <= U249_in;
    U5 <= U250_in;
    U6 <= U251_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X250_in;

    Y1 <= Y233_in;
    Y2 <= Y234_in;
    Y3 <= Y235_in;
    Y4 <= Y249_in;
    Y5 <= Y250_in;
    Y6 <= Y251_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11111010) begin // 251

    Y250_next <= Y_onebyoneout;
    X250_next <= X_onebyoneout;

    U1 <= U234_in;
    U2 <= U235_in;
    U3 <= U236_in;
    U4 <= U250_in;
    U5 <= U251_in;
    U6 <= U252_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X251_in;

    Y1 <= Y234_in;
    Y2 <= Y235_in;
    Y3 <= Y236_in;
    Y4 <= Y250_in;
    Y5 <= Y251_in;
    Y6 <= Y252_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11111011) begin // 252

    Y251_next <= Y_onebyoneout;
    X251_next <= X_onebyoneout;

    U1 <= U235_in;
    U2 <= U236_in;
    U3 <= U237_in;
    U4 <= U251_in;
    U5 <= U252_in;
    U6 <= U253_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X252_in;

    Y1 <= Y235_in;
    Y2 <= Y236_in;
    Y3 <= Y237_in;
    Y4 <= Y251_in;
    Y5 <= Y252_in;
    Y6 <= Y253_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11111100) begin // 253

    Y252_next <= Y_onebyoneout;
    X252_next <= X_onebyoneout;

    U1 <= U236_in;
    U2 <= U237_in;
    U3 <= U238_in;
    U4 <= U252_in;
    U5 <= U253_in;
    U6 <= U254_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X253_in;

    Y1 <= Y236_in;
    Y2 <= Y237_in;
    Y3 <= Y238_in;
    Y4 <= Y252_in;
    Y5 <= Y253_in;
    Y6 <= Y254_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11111101) begin // 254

    Y253_next <= Y_onebyoneout;
    X253_next <= X_onebyoneout;

    U1 <= U237_in;
    U2 <= U238_in;
    U3 <= U239_in;
    U4 <= U253_in;
    U5 <= U254_in;
    U6 <= U255_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X254_in;

    Y1 <= Y237_in;
    Y2 <= Y238_in;
    Y3 <= Y239_in;
    Y4 <= Y253_in;
    Y5 <= Y254_in;
    Y6 <= Y255_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11111110) begin // 255

    Y254_next <= Y_onebyoneout;
    X254_next <= X_onebyoneout;

    U1 <= U238_in;
    U2 <= U239_in;
    U3 <= U240_in;
    U4 <= U254_in;
    U5 <= U255_in;
    U6 <= U256_in;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X255_in;

    Y1 <= Y238_in;
    Y2 <= Y239_in;
    Y3 <= Y240_in;
    Y4 <= Y254_in;
    Y5 <= Y255_in;
    Y6 <= Y256_in;
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};


  end else if (counter == `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b11111111) begin // 256

    Y255_next <= Y_onebyoneout;
    X255_next <= X_onebyoneout;

    U1 <= U239_in;
    U2 <= U240_in;
    U3 <= `WIDTH'b0;
    U4 <= U255_in;
    U5 <= U256_in;
    U6 <= `WIDTH'b0;
    U7 <= `WIDTH'b0;
    U8 <= `WIDTH'b0;
    U9 <= `WIDTH'b0;

    X <= X256_in;

    Y1 <= Y239_in;
    Y2 <= Y240_in;
    Y3 <= {(2 * `WIDTH){1'b0}};
    Y4 <= Y255_in;
    Y5 <= Y256_in;
    Y6 <= {(2 * `WIDTH){1'b0}};
    Y7 <= {(2 * `WIDTH){1'b0}};
    Y8 <= {(2 * `WIDTH){1'b0}};
    Y9 <= {(2 * `WIDTH){1'b0}};

    end
  counter = counter + `COUNTER_WIDTH_SIXTEEN_BY_SIXTEEN'b1;
end

onebyone18mul u1(
.A1(A1[`WIDTH - 1:0]),
.A2(A2[`WIDTH - 1:0]),
.A3(A3[`WIDTH - 1:0]),
.A4(A4[`WIDTH - 1:0]),
.A5(A5[`WIDTH - 1:0]),
.A6(A6[`WIDTH - 1:0]),
.A7(A7[`WIDTH - 1:0]),
.A8(A8[`WIDTH - 1:0]),
.A9(A9[`WIDTH - 1:0]),

.B1(B1[`WIDTH - 1:0]),
.B2(B2[`WIDTH - 1:0]),
.B3(B3[`WIDTH - 1:0]),
.B4(B4[`WIDTH - 1:0]),
.B5(B5[`WIDTH - 1:0]),
.B6(B6[`WIDTH - 1:0]),
.B7(B7[`WIDTH - 1:0]),
.B8(B8[`WIDTH - 1:0]),
.B9(B9[`WIDTH - 1:0]),

.U1(U1[`WIDTH - 1:0]),
.U2(U2[`WIDTH - 1:0]),
.U3(U3[`WIDTH - 1:0]),
.U4(U4[`WIDTH - 1:0]),
.U5(U5[`WIDTH - 1:0]),
.U6(U6[`WIDTH - 1:0]),
.U7(U7[`WIDTH - 1:0]),
.U8(U8[`WIDTH - 1:0]),
.U9(U9[`WIDTH - 1:0]),

.Y1(Y1[2 * `WIDTH - 1:0]),
.Y2(Y2[2 * `WIDTH - 1:0]),
.Y3(Y3[2 * `WIDTH - 1:0]),
.Y4(Y4[2 * `WIDTH - 1:0]),
.Y5(Y5[2 * `WIDTH - 1:0]),
.Y6(Y6[2 * `WIDTH - 1:0]),
.Y7(Y7[2 * `WIDTH - 1:0]),
.Y8(Y8[2 * `WIDTH - 1:0]),
.Y9(Y9[2 * `WIDTH - 1:0]),

.I(I[`WIDTH - 1:0]),

.Xout(X_onebyoneout[2 * `WIDTH - 1:0]),
.Yout(Y_onebyoneout[2 * `WIDTH - 1:0]),
.X(X[2 * `WIDTH - 1:0])

);

endmodule
